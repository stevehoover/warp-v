`define RW_ZX(in, width) {{width-$width(in){1'b0}}, in}
