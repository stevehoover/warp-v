`ifndef SP_DEFAULT
`define SP_DEFAULT

// File included by SandPiper-generated code for the default project configuration.
`include "sandpiper.vh"


`endif  // SP_DEFAULT
