module clk_gate (output gated_clk, input free_clk, func_en, pwr_en, gating_override);

   assign gated_clk = free_clk;
endmodule
`ifndef SANDPIPER_VH
`define SANDPIPER_VH

`ifdef WHEN
   // Make sure user definition does not collide.
   !!!ERROR: WHEN macro already defined
`else
   `ifdef SP_PHYS
      // Phys compilation disabled X-injection.
      `define WHEN(valid_sig)
   `else
      // Inject X.
      `define WHEN(valid_sig) !valid_sig ? 'x :
   `endif
`endif

`endif


`define BOGUS_USE(ignore)
   
//include "sp_default.vh" //_\source warp-v_5-stage.tlv 5
//_\SV
   // Include WARP-V.
   // Included URL: "./warp-v.tlv"
//_\SV
module top(input logic clk, input logic reset, input logic [31:0] cyc_cnt, output logic passed, output logic failed);    /* verilator lint_save */ /* verilator lint_off UNOPTFLAT */ /* verilator lint_restore */  /* verilator lint_off WIDTH */ /* verilator lint_off UNOPTFLAT */
//_\source warp-v_5-stage.tlv 9
//`include "warp-v_5-stage_gen.sv"
// Generated by SandPiper(TM) 1.9-2018/02/11-beta from Redwood EDA.
// Redwood EDA does not claim intellectual property rights to this file and provides no warranty regarding its correctness or quality.


//`include "sandpiper_gen.vh"


genvar bank, instrs, mem, regs, src;


//
// Signals declared top-level.
//

// For |fetch/instr$Cnt.
logic [7:0] FETCH_Instr_Cnt_n2,
            FETCH_Instr_Cnt_n1;

// For |fetch/instr$GoodPathMask.
logic [1+1:0] FETCH_Instr_GoodPathMask_n1,
              FETCH_Instr_GoodPathMask_a0;

// For |fetch/instr$Pc.
logic [31:2] FETCH_Instr_Pc_n1,
             FETCH_Instr_Pc_a0;

// For |fetch/instr$ReachedEnd.
logic FETCH_Instr_ReachedEnd_n1,
      FETCH_Instr_ReachedEnd_a0;

// For |fetch/instr$Reg4Became45.
logic FETCH_Instr_Reg4Became45_n1,
      FETCH_Instr_Reg4Became45_a0;

// For |fetch/instr$RemainingCyclesWithinTimeUnit.
logic [30-1:0] FETCH_Instr_RemainingCyclesWithinTimeUnit_n1,
               FETCH_Instr_RemainingCyclesWithinTimeUnit_a0;

// For |fetch/instr$abort.
logic FETCH_Instr_abort_a0;

// For |fetch/instr$aborting_isa_trap.
logic FETCH_Instr_aborting_isa_trap_a0;

// For |fetch/instr$aborting_trap.
logic FETCH_Instr_aborting_trap_a0,
      FETCH_Instr_aborting_trap_a1;

// For |fetch/instr$add_sub_rslt.
logic [31:0] FETCH_Instr_add_sub_rslt_a0;

// For |fetch/instr$addi_rslt.
logic [31:0] FETCH_Instr_addi_rslt_a0;

// For |fetch/instr$addr.
logic [31:0] FETCH_Instr_addr_a0;

// For |fetch/instr$and_rslt.
logic [31:0] FETCH_Instr_and_rslt_a0;

// For |fetch/instr$andi_rslt.
logic [31:0] FETCH_Instr_andi_rslt_a0;

// For |fetch/instr$auipc_rslt.
logic [31:0] FETCH_Instr_auipc_rslt_a0;

// For |fetch/instr$branch.
logic FETCH_Instr_branch_a0;

// For |fetch/instr$branch_redir_pc.
logic [31:2] FETCH_Instr_branch_redir_pc_a0;

// For |fetch/instr$branch_target.
logic [31:2] FETCH_Instr_branch_target_a0;

// For |fetch/instr$commit.
logic FETCH_Instr_commit_a0,
      FETCH_Instr_commit_a1,
      FETCH_Instr_commit_a2,
      FETCH_Instr_commit_a3,
      FETCH_Instr_commit_a4,
      FETCH_Instr_commit_a5,
      FETCH_Instr_commit_a6;

// For |fetch/instr$conditional_branch.
logic FETCH_Instr_conditional_branch_a0;

// For |fetch/instr$csr_cycle.
logic [31:0] FETCH_Instr_csr_cycle_n1,
             FETCH_Instr_csr_cycle_a0;

// For |fetch/instr$csr_cycle_hw_wr.
logic FETCH_Instr_csr_cycle_hw_wr_a0;

// For |fetch/instr$csr_cycle_hw_wr_en_mask.
logic [31:0] FETCH_Instr_csr_cycle_hw_wr_en_mask_a0;

// For |fetch/instr$csr_cycle_hw_wr_mask.
logic FETCH_Instr_csr_cycle_hw_wr_mask_a0;

// For |fetch/instr$csr_cycle_hw_wr_value.
logic FETCH_Instr_csr_cycle_hw_wr_value_a0;

// For |fetch/instr$csr_cycle_masked_wr_value.
logic [31:0] FETCH_Instr_csr_cycle_masked_wr_value_a0;

// For |fetch/instr$csr_cycleh.
logic [31:0] FETCH_Instr_csr_cycleh_n1,
             FETCH_Instr_csr_cycleh_a0;

// For |fetch/instr$csr_cycleh_hw_wr.
logic FETCH_Instr_csr_cycleh_hw_wr_a0;

// For |fetch/instr$csr_cycleh_hw_wr_en_mask.
logic [31:0] FETCH_Instr_csr_cycleh_hw_wr_en_mask_a0;

// For |fetch/instr$csr_cycleh_hw_wr_mask.
logic FETCH_Instr_csr_cycleh_hw_wr_mask_a0;

// For |fetch/instr$csr_cycleh_hw_wr_value.
logic FETCH_Instr_csr_cycleh_hw_wr_value_a0;

// For |fetch/instr$csr_cycleh_masked_wr_value.
logic [31:0] FETCH_Instr_csr_cycleh_masked_wr_value_a0;

// For |fetch/instr$csr_instret.
logic [31:0] FETCH_Instr_csr_instret_n1,
             FETCH_Instr_csr_instret_a0;

// For |fetch/instr$csr_instret_hw_wr.
logic FETCH_Instr_csr_instret_hw_wr_a0;

// For |fetch/instr$csr_instret_hw_wr_en_mask.
logic [31:0] FETCH_Instr_csr_instret_hw_wr_en_mask_a0;

// For |fetch/instr$csr_instret_hw_wr_mask.
logic FETCH_Instr_csr_instret_hw_wr_mask_a0;

// For |fetch/instr$csr_instret_hw_wr_value.
logic FETCH_Instr_csr_instret_hw_wr_value_a0;

// For |fetch/instr$csr_instret_masked_wr_value.
logic [31:0] FETCH_Instr_csr_instret_masked_wr_value_a0;

// For |fetch/instr$csr_instreth.
logic [31:0] FETCH_Instr_csr_instreth_n1,
             FETCH_Instr_csr_instreth_a0;

// For |fetch/instr$csr_instreth_hw_wr.
logic FETCH_Instr_csr_instreth_hw_wr_a0;

// For |fetch/instr$csr_instreth_hw_wr_en_mask.
logic [31:0] FETCH_Instr_csr_instreth_hw_wr_en_mask_a0;

// For |fetch/instr$csr_instreth_hw_wr_mask.
logic FETCH_Instr_csr_instreth_hw_wr_mask_a0;

// For |fetch/instr$csr_instreth_hw_wr_value.
logic FETCH_Instr_csr_instreth_hw_wr_value_a0;

// For |fetch/instr$csr_instreth_masked_wr_value.
logic [31:0] FETCH_Instr_csr_instreth_masked_wr_value_a0;

// For |fetch/instr$csr_time.
logic [31:0] FETCH_Instr_csr_time_n1,
             FETCH_Instr_csr_time_a0;

// For |fetch/instr$csr_time_hw_wr.
logic FETCH_Instr_csr_time_hw_wr_a0;

// For |fetch/instr$csr_time_hw_wr_en_mask.
logic [31:0] FETCH_Instr_csr_time_hw_wr_en_mask_a0;

// For |fetch/instr$csr_time_hw_wr_mask.
logic FETCH_Instr_csr_time_hw_wr_mask_a0;

// For |fetch/instr$csr_time_hw_wr_value.
logic FETCH_Instr_csr_time_hw_wr_value_a0;

// For |fetch/instr$csr_time_masked_wr_value.
logic [31:0] FETCH_Instr_csr_time_masked_wr_value_a0;

// For |fetch/instr$csr_timeh.
logic [31:0] FETCH_Instr_csr_timeh_n1,
             FETCH_Instr_csr_timeh_a0;

// For |fetch/instr$csr_timeh_hw_wr.
logic FETCH_Instr_csr_timeh_hw_wr_a0;

// For |fetch/instr$csr_timeh_hw_wr_en_mask.
logic [31:0] FETCH_Instr_csr_timeh_hw_wr_en_mask_a0;

// For |fetch/instr$csr_timeh_hw_wr_mask.
logic FETCH_Instr_csr_timeh_hw_wr_mask_a0;

// For |fetch/instr$csr_timeh_hw_wr_value.
logic FETCH_Instr_csr_timeh_hw_wr_value_a0;

// For |fetch/instr$csr_timeh_masked_wr_value.
logic [31:0] FETCH_Instr_csr_timeh_masked_wr_value_a0;

// For |fetch/instr$csr_trap.
logic FETCH_Instr_csr_trap_a0;

// For |fetch/instr$csrrc_rslt.
logic [31:0] FETCH_Instr_csrrc_rslt_a0;

// For |fetch/instr$csrrci_rslt.
logic [31:0] FETCH_Instr_csrrci_rslt_a0;

// For |fetch/instr$csrrs_rslt.
logic [31:0] FETCH_Instr_csrrs_rslt_a0;

// For |fetch/instr$csrrsi_rslt.
logic [31:0] FETCH_Instr_csrrsi_rslt_a0;

// For |fetch/instr$csrrw_rslt.
logic [31:0] FETCH_Instr_csrrw_rslt_a0;

// For |fetch/instr$csrrwi_rslt.
logic [31:0] FETCH_Instr_csrrwi_rslt_a0;

// For |fetch/instr$dest_pending.
logic FETCH_Instr_dest_pending_a0;

// For |fetch/instr$dest_reg.
logic [4:0] FETCH_Instr_dest_reg_a0;

// For |fetch/instr$dest_reg_valid.
logic FETCH_Instr_dest_reg_valid_a0;

// For |fetch/instr$equal.
logic FETCH_Instr_equal_a0;

// For |fetch/instr$fetch.
logic FETCH_Instr_fetch_a0;

// For |fetch/instr$full_csr_cycle_hw_wr_value.
logic [63:0] FETCH_Instr_full_csr_cycle_hw_wr_value_a0;

// For |fetch/instr$full_csr_instret_hw_wr_value.
logic [63:0] FETCH_Instr_full_csr_instret_hw_wr_value_a0;

// For |fetch/instr$full_csr_time_hw_wr_value.
logic [63:0] FETCH_Instr_full_csr_time_hw_wr_value_a0;

// For |fetch/instr$illegal.
logic FETCH_Instr_illegal_a0,
      FETCH_Instr_illegal_a1,
      FETCH_Instr_illegal_a2,
      FETCH_Instr_illegal_a3,
      FETCH_Instr_illegal_a4,
      FETCH_Instr_illegal_a5,
      FETCH_Instr_illegal_a6;

// For |fetch/instr$indirect_jump.
logic FETCH_Instr_indirect_jump_a0;

// For |fetch/instr$indirect_jump_full_target.
logic [31:0] FETCH_Instr_indirect_jump_full_target_a0;

// For |fetch/instr$indirect_jump_target.
logic [31:2] FETCH_Instr_indirect_jump_target_a0;

// For |fetch/instr$is___type.
logic FETCH_Instr_is___type_a0;

// For |fetch/instr$is_add_sub_instr.
logic FETCH_Instr_is_add_sub_instr_a0;

// For |fetch/instr$is_addi_instr.
logic FETCH_Instr_is_addi_instr_a0;

// For |fetch/instr$is_and_instr.
logic FETCH_Instr_is_and_instr_a0;

// For |fetch/instr$is_andi_instr.
logic FETCH_Instr_is_andi_instr_a0;

// For |fetch/instr$is_auipc_instr.
logic FETCH_Instr_is_auipc_instr_a0;

// For |fetch/instr$is_b_type.
logic FETCH_Instr_is_b_type_a0;

// For |fetch/instr$is_beq_instr.
logic FETCH_Instr_is_beq_instr_a0;

// For |fetch/instr$is_bge_instr.
logic FETCH_Instr_is_bge_instr_a0;

// For |fetch/instr$is_bgeu_instr.
logic FETCH_Instr_is_bgeu_instr_a0;

// For |fetch/instr$is_blt_instr.
logic FETCH_Instr_is_blt_instr_a0;

// For |fetch/instr$is_bltu_instr.
logic FETCH_Instr_is_bltu_instr_a0;

// For |fetch/instr$is_bne_instr.
logic FETCH_Instr_is_bne_instr_a0;

// For |fetch/instr$is_csr_cycle.
logic FETCH_Instr_is_csr_cycle_a0;

// For |fetch/instr$is_csr_cycleh.
logic FETCH_Instr_is_csr_cycleh_a0;

// For |fetch/instr$is_csr_instr.
logic FETCH_Instr_is_csr_instr_a0;

// For |fetch/instr$is_csr_instret.
logic FETCH_Instr_is_csr_instret_a0;

// For |fetch/instr$is_csr_instreth.
logic FETCH_Instr_is_csr_instreth_a0;

// For |fetch/instr$is_csr_time.
logic FETCH_Instr_is_csr_time_a0;

// For |fetch/instr$is_csr_timeh.
logic FETCH_Instr_is_csr_timeh_a0;

// For |fetch/instr$is_csrrc_instr.
logic FETCH_Instr_is_csrrc_instr_a0;

// For |fetch/instr$is_csrrci_instr.
logic FETCH_Instr_is_csrrci_instr_a0;

// For |fetch/instr$is_csrrs_instr.
logic FETCH_Instr_is_csrrs_instr_a0;

// For |fetch/instr$is_csrrsi_instr.
logic FETCH_Instr_is_csrrsi_instr_a0;

// For |fetch/instr$is_csrrw_instr.
logic FETCH_Instr_is_csrrw_instr_a0;

// For |fetch/instr$is_csrrwi_instr.
logic FETCH_Instr_is_csrrwi_instr_a0;

// For |fetch/instr$is_dest_condition.
logic FETCH_Instr_is_dest_condition_a0;

// For |fetch/instr$is_i_type.
logic FETCH_Instr_is_i_type_a0;

// For |fetch/instr$is_j_type.
logic FETCH_Instr_is_j_type_a0;

// For |fetch/instr$is_jal_instr.
logic FETCH_Instr_is_jal_instr_a0;

// For |fetch/instr$is_jalr_instr.
logic FETCH_Instr_is_jalr_instr_a0;

// For |fetch/instr$is_lb_instr.
logic FETCH_Instr_is_lb_instr_a0;

// For |fetch/instr$is_lbu_instr.
logic FETCH_Instr_is_lbu_instr_a0;

// For |fetch/instr$is_lh_instr.
logic FETCH_Instr_is_lh_instr_a0;

// For |fetch/instr$is_lhu_instr.
logic FETCH_Instr_is_lhu_instr_a0;

// For |fetch/instr$is_lui_instr.
logic FETCH_Instr_is_lui_instr_a0;

// For |fetch/instr$is_lw_instr.
logic FETCH_Instr_is_lw_instr_a0;

// For |fetch/instr$is_or_instr.
logic FETCH_Instr_is_or_instr_a0;

// For |fetch/instr$is_ori_instr.
logic FETCH_Instr_is_ori_instr_a0;

// For |fetch/instr$is_r4_type.
logic FETCH_Instr_is_r4_type_a0;

// For |fetch/instr$is_r_type.
logic FETCH_Instr_is_r_type_a0;

// For |fetch/instr$is_ri_type.
logic FETCH_Instr_is_ri_type_a0;

// For |fetch/instr$is_s_type.
logic FETCH_Instr_is_s_type_a0;

// For |fetch/instr$is_sb_instr.
logic FETCH_Instr_is_sb_instr_a0;

// For |fetch/instr$is_sh_instr.
logic FETCH_Instr_is_sh_instr_a0;

// For |fetch/instr$is_sll_instr.
logic FETCH_Instr_is_sll_instr_a0;

// For |fetch/instr$is_slli_instr.
logic FETCH_Instr_is_slli_instr_a0;

// For |fetch/instr$is_slt_instr.
logic FETCH_Instr_is_slt_instr_a0;

// For |fetch/instr$is_slti_instr.
logic FETCH_Instr_is_slti_instr_a0;

// For |fetch/instr$is_sltiu_instr.
logic FETCH_Instr_is_sltiu_instr_a0;

// For |fetch/instr$is_sltu_instr.
logic FETCH_Instr_is_sltu_instr_a0;

// For |fetch/instr$is_srl_sra_instr.
logic FETCH_Instr_is_srl_sra_instr_a0;

// For |fetch/instr$is_srli_srai_instr.
logic FETCH_Instr_is_srli_srai_instr_a0;

// For |fetch/instr$is_sw_instr.
logic FETCH_Instr_is_sw_instr_a0;

// For |fetch/instr$is_u_type.
logic FETCH_Instr_is_u_type_a0;

// For |fetch/instr$is_xor_instr.
logic FETCH_Instr_is_xor_instr_a0;

// For |fetch/instr$is_xori_instr.
logic FETCH_Instr_is_xori_instr_a0;

// For |fetch/instr$jal_rslt.
logic [31:0] FETCH_Instr_jal_rslt_a0;

// For |fetch/instr$jalr_rslt.
logic [31:0] FETCH_Instr_jalr_rslt_a0;

// For |fetch/instr$jump.
logic FETCH_Instr_jump_a0;

// For |fetch/instr$jump_target.
logic [31:2] FETCH_Instr_jump_target_a0;

// For |fetch/instr$lb_rslt.
logic [31:0] FETCH_Instr_lb_rslt_a0;

// For |fetch/instr$lbu_rslt.
logic [31:0] FETCH_Instr_lbu_rslt_a0;

// For |fetch/instr$ld.
logic FETCH_Instr_ld_a0;

// For |fetch/instr$ld_st.
logic FETCH_Instr_ld_st_a0;

// For |fetch/instr$ld_st_cond.
logic FETCH_Instr_ld_st_cond_a0;

// For |fetch/instr$ld_st_half.
logic FETCH_Instr_ld_st_half_a0;

// For |fetch/instr$ld_st_word.
logic FETCH_Instr_ld_st_word_a0;

// For |fetch/instr$ld_value.
logic [31:0] FETCH_Instr_ld_value_a0;

// For |fetch/instr$lh_rslt.
logic [31:0] FETCH_Instr_lh_rslt_a0;

// For |fetch/instr$lhu_rslt.
logic [31:0] FETCH_Instr_lhu_rslt_a0;

// For |fetch/instr$lui_rslt.
logic [31:0] FETCH_Instr_lui_rslt_a0;

// For |fetch/instr$lw_rslt.
logic [31:0] FETCH_Instr_lw_rslt_a0;

// For |fetch/instr$masked_csr_wr_value.
logic [31:0] FETCH_Instr_masked_csr_wr_value_a0;

// For |fetch/instr$misaligned_indirect_jump_target.
logic FETCH_Instr_misaligned_indirect_jump_target_a0;

// For |fetch/instr$misaligned_jump_target.
logic FETCH_Instr_misaligned_jump_target_a0;

// For |fetch/instr$misaligned_pc.
logic FETCH_Instr_misaligned_pc_a0;

// For |fetch/instr$mispred_branch.
logic FETCH_Instr_mispred_branch_a0;

// For |fetch/instr$mnemonic.
logic [10*8-1:0] FETCH_Instr_mnemonic_a0;

// For |fetch/instr$next_good_path_mask.
logic [1+1:0] FETCH_Instr_next_good_path_mask_a0;

// For |fetch/instr$non_aborting_isa_trap.
logic FETCH_Instr_non_aborting_isa_trap_a0;

// For |fetch/instr$non_aborting_trap.
logic FETCH_Instr_non_aborting_trap_a0,
      FETCH_Instr_non_aborting_trap_a1;

// For |fetch/instr$or_rslt.
logic [31:0] FETCH_Instr_or_rslt_a0;

// For |fetch/instr$ori_rslt.
logic [31:0] FETCH_Instr_ori_rslt_a0;

// For |fetch/instr$pred_taken.
logic FETCH_Instr_pred_taken_a0;

// For |fetch/instr$raw.
logic [31:0] FETCH_Instr_raw_a0;

// For |fetch/instr$raw_aq.
logic FETCH_Instr_raw_aq_a0;

// For |fetch/instr$raw_b_imm.
logic [31:0] FETCH_Instr_raw_b_imm_a0;

// For |fetch/instr$raw_funct3.
logic [2:0] FETCH_Instr_raw_funct3_a0;

// For |fetch/instr$raw_funct7.
logic [6:0] FETCH_Instr_raw_funct7_a0;

// For |fetch/instr$raw_i_imm.
logic [31:0] FETCH_Instr_raw_i_imm_a0;

// For |fetch/instr$raw_j_imm.
logic [31:0] FETCH_Instr_raw_j_imm_a0;

// For |fetch/instr$raw_op2.
logic [1:0] FETCH_Instr_raw_op2_a0;

// For |fetch/instr$raw_op5.
logic [4:0] FETCH_Instr_raw_op5_a0;

// For |fetch/instr$raw_rd.
logic [4:0] FETCH_Instr_raw_rd_a0;

// For |fetch/instr$raw_rl.
logic FETCH_Instr_raw_rl_a0;

// For |fetch/instr$raw_rm.
logic [2:0] FETCH_Instr_raw_rm_a0;

// For |fetch/instr$raw_rs1.
logic [4:0] FETCH_Instr_raw_rs1_a0;

// For |fetch/instr$raw_rs2.
logic [4:0] FETCH_Instr_raw_rs2_a0;

// For |fetch/instr$raw_rs3.
logic [4:0] FETCH_Instr_raw_rs3_a0;

// For |fetch/instr$raw_s_imm.
logic [31:0] FETCH_Instr_raw_s_imm_a0;

// For |fetch/instr$raw_shamt.
logic [6:0] FETCH_Instr_raw_shamt_a0;

// For |fetch/instr$raw_u_imm.
logic [31:0] FETCH_Instr_raw_u_imm_a0;

// For |fetch/instr$reg_wr_pending.
logic FETCH_Instr_reg_wr_pending_a0;

// For |fetch/instr$reg_write.
logic FETCH_Instr_reg_write_a0;

// For |fetch/instr$replay.
logic FETCH_Instr_replay_a0,
      FETCH_Instr_replay_a1;

// For |fetch/instr$reset.
logic FETCH_Instr_reset_n1,
      FETCH_Instr_reset_a0,
      FETCH_Instr_reset_a1,
      FETCH_Instr_reset_a2,
      FETCH_Instr_reset_a3;

// For |fetch/instr$returning_ld.
logic FETCH_Instr_returning_ld_a0,
      FETCH_Instr_returning_ld_a1;

// For |fetch/instr$rslt.
logic [31:0] FETCH_Instr_rslt_a0;

// For |fetch/instr$sll_rslt.
logic [31:0] FETCH_Instr_sll_rslt_a0;

// For |fetch/instr$slli_rslt.
logic [31:0] FETCH_Instr_slli_rslt_a0;

// For |fetch/instr$slt_rslt.
logic [31:0] FETCH_Instr_slt_rslt_a0;

// For |fetch/instr$slti_rslt.
logic [31:0] FETCH_Instr_slti_rslt_a0;

// For |fetch/instr$sltiu_rslt.
logic [31:0] FETCH_Instr_sltiu_rslt_a0;

// For |fetch/instr$sltu_rslt.
logic [31:0] FETCH_Instr_sltu_rslt_a0;

// For |fetch/instr$spec_ld.
logic FETCH_Instr_spec_ld_a0;

// For |fetch/instr$sra_intermediate_rslt.
logic [31:0] FETCH_Instr_sra_intermediate_rslt_a0;

// For |fetch/instr$srai_intermediate_rslt.
logic [31:0] FETCH_Instr_srai_intermediate_rslt_a0;

// For |fetch/instr$srl_intermediate_rslt.
logic [31:0] FETCH_Instr_srl_intermediate_rslt_a0;

// For |fetch/instr$srl_sra_rslt.
logic [31:0] FETCH_Instr_srl_sra_rslt_a0;

// For |fetch/instr$srli_intermediate_rslt.
logic [31:0] FETCH_Instr_srli_intermediate_rslt_a0;

// For |fetch/instr$srli_srai_rslt.
logic [31:0] FETCH_Instr_srli_srai_rslt_a0;

// For |fetch/instr$st.
logic FETCH_Instr_st_a0;

// For |fetch/instr$st_cond.
logic FETCH_Instr_st_cond_a0;

// For |fetch/instr$st_mask.
logic [3:0] FETCH_Instr_st_mask_a0;

// For |fetch/instr$st_reg_value.
logic [31:0] FETCH_Instr_st_reg_value_a0;

// For |fetch/instr$st_value.
logic [31:0] FETCH_Instr_st_value_a0;

// For |fetch/instr$taken.
logic FETCH_Instr_taken_a0;

// For |fetch/instr$time_unit_expires.
logic FETCH_Instr_time_unit_expires_a0;

// For |fetch/instr$trap_target.
logic [31:2] FETCH_Instr_trap_target_a0,
             FETCH_Instr_trap_target_a1;

// For |fetch/instr$unnatural_addr_trap.
logic FETCH_Instr_unnatural_addr_trap_a0;

// For |fetch/instr$upd_csr_cycle.
logic [31:0] FETCH_Instr_upd_csr_cycle_a0;

// For |fetch/instr$upd_csr_cycleh.
logic [31:0] FETCH_Instr_upd_csr_cycleh_a0;

// For |fetch/instr$upd_csr_instret.
logic [31:0] FETCH_Instr_upd_csr_instret_a0;

// For |fetch/instr$upd_csr_instreth.
logic [31:0] FETCH_Instr_upd_csr_instreth_a0;

// For |fetch/instr$upd_csr_time.
logic [31:0] FETCH_Instr_upd_csr_time_a0;

// For |fetch/instr$upd_csr_timeh.
logic [31:0] FETCH_Instr_upd_csr_timeh_a0;

// For |fetch/instr$valid_csr.
logic FETCH_Instr_valid_csr_a0;

// For |fetch/instr$valid_decode.
logic FETCH_Instr_valid_decode_a0,
      FETCH_Instr_valid_decode_a1,
      FETCH_Instr_valid_decode_a2,
      FETCH_Instr_valid_decode_a3,
      FETCH_Instr_valid_decode_a4,
      FETCH_Instr_valid_decode_a5;

// For |fetch/instr$valid_decode_branch.
logic FETCH_Instr_valid_decode_branch_a0;

// For |fetch/instr$valid_dest_reg_valid.
logic FETCH_Instr_valid_dest_reg_valid_a0;

// For |fetch/instr$valid_exe.
logic FETCH_Instr_valid_exe_a0;

// For |fetch/instr$valid_ld.
logic FETCH_Instr_valid_ld_a0;

// For |fetch/instr$valid_st.
logic FETCH_Instr_valid_st_a0;

// For |fetch/instr$xor_rslt.
logic [31:0] FETCH_Instr_xor_rslt_a0;

// For |fetch/instr$xori_rslt.
logic [31:0] FETCH_Instr_xori_rslt_a0;

// For |fetch/instr/original_ld$addr.
logic [1:0] FETCH_Instr_OriginalLd_addr_a0;

// For |fetch/instr/original_ld$dest_reg.
logic [4:0] FETCH_Instr_OriginalLd_dest_reg_a0;

// For |fetch/instr/original_ld$ld_mask.
logic [3:0] FETCH_Instr_OriginalLd_ld_mask_a0;

// For |fetch/instr/original_ld$ld_rslt.
logic [31:0] FETCH_Instr_OriginalLd_ld_rslt_a0;

// For |fetch/instr/original_ld$ld_st_half.
logic FETCH_Instr_OriginalLd_ld_st_half_a0;

// For |fetch/instr/original_ld$ld_st_word.
logic FETCH_Instr_OriginalLd_ld_st_word_a0;

// For |fetch/instr/original_ld$ld_value.
logic [31:0] FETCH_Instr_OriginalLd_ld_value_a0;

// For |fetch/instr/original_ld$raw_funct3.
logic [2:2] FETCH_Instr_OriginalLd_raw_funct3_a0;

// For |fetch/instr/original_ld$sign_bit.
logic FETCH_Instr_OriginalLd_sign_bit_a0;

// For |fetch/instr/regs$pending.
logic FETCH_Instr_Regs_pending_n1 [31:1],
      FETCH_Instr_Regs_pending_a0 [31:1];

// For |fetch/instr/regs$value.
logic [31:0] FETCH_Instr_Regs_value_a0 [31:1];

// For |fetch/instr/src$replay.
logic [2:1] FETCH_Instr_Src_replay_a0;

// For |fetch/instrs$instr.
logic [31:0] FETCH_Instrs_instr_a0 [11:0];

// For |mem/data$addr.
logic [1:0] MEM_Data_addr_a0,
            MEM_Data_addr_a1;

// For |mem/data$dest_reg.
logic [4:0] MEM_Data_dest_reg_a0,
            MEM_Data_dest_reg_a1;

// For |mem/data$ld_st_half.
logic MEM_Data_ld_st_half_a0,
      MEM_Data_ld_st_half_a1;

// For |mem/data$ld_st_word.
logic MEM_Data_ld_st_word_a0,
      MEM_Data_ld_st_word_a1;

// For |mem/data$ld_value.
logic [31:0] MEM_Data_ld_value_a0,
             MEM_Data_ld_value_a1;

// For |mem/data$raw_funct3.
logic [2:2] MEM_Data_raw_funct3_a0,
            MEM_Data_raw_funct3_a1;

// For |mem/data$valid_ld.
logic MEM_Data_valid_ld_a0,
      MEM_Data_valid_ld_a1;


//
// Scope: |fetch
//

//
// Scope: |fetch/instr
//

// Clock signals.
logic clkP_FETCH_Instr_valid_decode_a1 ;
logic clkP_FETCH_Instr_valid_decode_a2 ;
logic clkP_FETCH_Instr_valid_decode_a3 ;
logic clkP_FETCH_Instr_valid_decode_a4 ;
logic clkP_FETCH_Instr_valid_decode_a5 ;
logic clkP_FETCH_Instr_valid_decode_a6 ;


generate


   //
   // Scope: |fetch
   //


      //
      // Scope: /instr
      //

         // For $Cnt.
         always_ff @(posedge clk) FETCH_Instr_Cnt_n1[7:0] <= FETCH_Instr_Cnt_n2[7:0];

         // For $GoodPathMask.
         always_ff @(posedge clk) FETCH_Instr_GoodPathMask_a0[1+1:0] <= FETCH_Instr_GoodPathMask_n1[1+1:0];

         // For $Pc.
         always_ff @(posedge clk) FETCH_Instr_Pc_a0[31:2] <= FETCH_Instr_Pc_n1[31:2];

         // For $ReachedEnd.
         always_ff @(posedge clk) FETCH_Instr_ReachedEnd_a0 <= FETCH_Instr_ReachedEnd_n1;

         // For $Reg4Became45.
         always_ff @(posedge clk) FETCH_Instr_Reg4Became45_a0 <= FETCH_Instr_Reg4Became45_n1;

         // For $RemainingCyclesWithinTimeUnit.
         always_ff @(posedge clk) FETCH_Instr_RemainingCyclesWithinTimeUnit_a0[30-1:0] <= FETCH_Instr_RemainingCyclesWithinTimeUnit_n1[30-1:0];

         // For $aborting_trap.
         always_ff @(posedge clk) FETCH_Instr_aborting_trap_a1 <= FETCH_Instr_aborting_trap_a0;

         // For $commit.
         always_ff @(posedge clk) FETCH_Instr_commit_a1 <= FETCH_Instr_commit_a0;
         always_ff @(posedge clk) FETCH_Instr_commit_a2 <= FETCH_Instr_commit_a1;
         always_ff @(posedge clk) FETCH_Instr_commit_a3 <= FETCH_Instr_commit_a2;
         always_ff @(posedge clk) FETCH_Instr_commit_a4 <= FETCH_Instr_commit_a3;
         always_ff @(posedge clk) FETCH_Instr_commit_a5 <= FETCH_Instr_commit_a4;
         always_ff @(posedge clk) FETCH_Instr_commit_a6 <= FETCH_Instr_commit_a5;

         // For $csr_cycle.
         always_ff @(posedge clk) FETCH_Instr_csr_cycle_a0[31:0] <= FETCH_Instr_csr_cycle_n1[31:0];

         // For $csr_cycleh.
         always_ff @(posedge clk) FETCH_Instr_csr_cycleh_a0[31:0] <= FETCH_Instr_csr_cycleh_n1[31:0];

         // For $csr_instret.
         always_ff @(posedge clk) FETCH_Instr_csr_instret_a0[31:0] <= FETCH_Instr_csr_instret_n1[31:0];

         // For $csr_instreth.
         always_ff @(posedge clk) FETCH_Instr_csr_instreth_a0[31:0] <= FETCH_Instr_csr_instreth_n1[31:0];

         // For $csr_time.
         always_ff @(posedge clk) FETCH_Instr_csr_time_a0[31:0] <= FETCH_Instr_csr_time_n1[31:0];

         // For $csr_timeh.
         always_ff @(posedge clk) FETCH_Instr_csr_timeh_a0[31:0] <= FETCH_Instr_csr_timeh_n1[31:0];

         // For $illegal.
         always_ff @(posedge clkP_FETCH_Instr_valid_decode_a1) FETCH_Instr_illegal_a1 <= FETCH_Instr_illegal_a0;
         always_ff @(posedge clkP_FETCH_Instr_valid_decode_a2) FETCH_Instr_illegal_a2 <= FETCH_Instr_illegal_a1;
         always_ff @(posedge clkP_FETCH_Instr_valid_decode_a3) FETCH_Instr_illegal_a3 <= FETCH_Instr_illegal_a2;
         always_ff @(posedge clkP_FETCH_Instr_valid_decode_a4) FETCH_Instr_illegal_a4 <= FETCH_Instr_illegal_a3;
         always_ff @(posedge clkP_FETCH_Instr_valid_decode_a5) FETCH_Instr_illegal_a5 <= FETCH_Instr_illegal_a4;
         always_ff @(posedge clkP_FETCH_Instr_valid_decode_a6) FETCH_Instr_illegal_a6 <= FETCH_Instr_illegal_a5;

         // For $non_aborting_trap.
         always_ff @(posedge clk) FETCH_Instr_non_aborting_trap_a1 <= FETCH_Instr_non_aborting_trap_a0;

         // For $replay.
         always_ff @(posedge clk) FETCH_Instr_replay_a1 <= FETCH_Instr_replay_a0;

         // For $reset.
         always_ff @(posedge clk) FETCH_Instr_reset_a0 <= FETCH_Instr_reset_n1;
         always_ff @(posedge clk) FETCH_Instr_reset_a1 <= FETCH_Instr_reset_a0;
         always_ff @(posedge clk) FETCH_Instr_reset_a2 <= FETCH_Instr_reset_a1;
         always_ff @(posedge clk) FETCH_Instr_reset_a3 <= FETCH_Instr_reset_a2;

         // For $returning_ld.
         always_ff @(posedge clk) FETCH_Instr_returning_ld_a1 <= FETCH_Instr_returning_ld_a0;

         // For $trap_target.
         always_ff @(posedge clk) FETCH_Instr_trap_target_a1[31:2] <= FETCH_Instr_trap_target_a0[31:2];

         // For $valid_decode.
         always_ff @(posedge clk) FETCH_Instr_valid_decode_a1 <= FETCH_Instr_valid_decode_a0;
         always_ff @(posedge clk) FETCH_Instr_valid_decode_a2 <= FETCH_Instr_valid_decode_a1;
         always_ff @(posedge clk) FETCH_Instr_valid_decode_a3 <= FETCH_Instr_valid_decode_a2;
         always_ff @(posedge clk) FETCH_Instr_valid_decode_a4 <= FETCH_Instr_valid_decode_a3;
         always_ff @(posedge clk) FETCH_Instr_valid_decode_a5 <= FETCH_Instr_valid_decode_a4;


         //
         // Scope: /regs[31:1]
         //
         for (regs = 1; regs <= 31; regs++) begin : L1gen_FETCH_Instr_Regs
            // For $pending.
            always_ff @(posedge clk) FETCH_Instr_Regs_pending_a0[regs] <= FETCH_Instr_Regs_pending_n1[regs];

         end



   //
   // Scope: |mem
   //


      //
      // Scope: /data
      //

         // For $addr.
         always_ff @(posedge clk) MEM_Data_addr_a1[1:0] <= MEM_Data_addr_a0[1:0];

         // For $dest_reg.
         always_ff @(posedge clk) MEM_Data_dest_reg_a1[4:0] <= MEM_Data_dest_reg_a0[4:0];

         // For $ld_st_half.
         always_ff @(posedge clk) MEM_Data_ld_st_half_a1 <= MEM_Data_ld_st_half_a0;

         // For $ld_st_word.
         always_ff @(posedge clk) MEM_Data_ld_st_word_a1 <= MEM_Data_ld_st_word_a0;

         // For $ld_value.
         always_ff @(posedge clk) MEM_Data_ld_value_a1[31:0] <= MEM_Data_ld_value_a0[31:0];

         // For $raw_funct3.
         always_ff @(posedge clk) MEM_Data_raw_funct3_a1[2] <= MEM_Data_raw_funct3_a0[2];

         // For $valid_ld.
         always_ff @(posedge clk) MEM_Data_valid_ld_a1 <= MEM_Data_valid_ld_a0;


         //
         // Scope: /src[2:1]
         //
         for (src = 1; src <= 2; src++) begin : L1gen_MEM_Data_Src
            // For $dummy.
            always_ff @(posedge clk) L1_MEM_Data_Src[src].L1_dummy_a1 <= L1_MEM_Data_Src[src].L1_dummy_a0;

         end




endgenerate



//
// Gated clocks.
//

generate



   //
   // Scope: |fetch
   //


      //
      // Scope: /instr
      //

         clk_gate gen_clkP_FETCH_Instr_valid_decode_a1(clkP_FETCH_Instr_valid_decode_a1, clk, 1'b1, FETCH_Instr_valid_decode_a0, 1'b0);
         clk_gate gen_clkP_FETCH_Instr_valid_decode_a2(clkP_FETCH_Instr_valid_decode_a2, clk, 1'b1, FETCH_Instr_valid_decode_a1, 1'b0);
         clk_gate gen_clkP_FETCH_Instr_valid_decode_a3(clkP_FETCH_Instr_valid_decode_a3, clk, 1'b1, FETCH_Instr_valid_decode_a2, 1'b0);
         clk_gate gen_clkP_FETCH_Instr_valid_decode_a4(clkP_FETCH_Instr_valid_decode_a4, clk, 1'b1, FETCH_Instr_valid_decode_a3, 1'b0);
         clk_gate gen_clkP_FETCH_Instr_valid_decode_a5(clkP_FETCH_Instr_valid_decode_a5, clk, 1'b1, FETCH_Instr_valid_decode_a4, 1'b0);
         clk_gate gen_clkP_FETCH_Instr_valid_decode_a6(clkP_FETCH_Instr_valid_decode_a6, clk, 1'b1, FETCH_Instr_valid_decode_a5, 1'b0);




endgenerate
generate //_\TLV
   //_\source ./warpv.tlv 1764   // Instantiated from warp-v_5-stage.tlv, 11 as: m4+cpu()
      
      // Generated logic
      //_\source <builtin> 1   // Instantiated from warp-v_5-stage.tlv, 1767 as: m4+indirect(M4_isa['_gen'])
         //_\source ./warpv.tlv 1142   // Instantiated from built-in definition.
         
            
            // v---------------------
            // Instruction characterization
         
            // M4 ugliness for instruction characterization.
            
            // For each opcode[6:2]
            // (User ISA Manual 2.2, Table 19.1)
            // Associate opcode[6:2] ([1:0] are 2'b11) with mnemonic and instruction type.
            // Instruction type is not in the table, but there seems to be a single instruction type for each of these,
            // so that is mapped here as well.
            // op5(bits, type, mnemonic)
            /*SV_plus*/
               localparam [4:0] OP5_LOAD = 5'b00000;
               localparam [4:0] OP5_LOAD_FP = 5'b00001;
               localparam [4:0] OP5_CUSTOM_0 = 5'b00010;
               localparam [4:0] OP5_MISC_MEM = 5'b00011;
               localparam [4:0] OP5_OP_IMM = 5'b00100;
               localparam [4:0] OP5_AUIPC = 5'b00101;
               localparam [4:0] OP5_OP_IMM_32 = 5'b00110;
               localparam [4:0] OP5_48B1 = 5'b00111;
               localparam [4:0] OP5_STORE = 5'b01000;
               localparam [4:0] OP5_STORE_FP = 5'b01001;
               localparam [4:0] OP5_CUSTOM_1 = 5'b01010;
               localparam [4:0] OP5_AMO = 5'b01011;  // (R-type, but rs2 = const for some, based on funct7 which doesn't exist for I-type?? R-type w/ ignored R2?)
               localparam [4:0] OP5_OP = 5'b01100;
               localparam [4:0] OP5_LUI = 5'b01101;
               localparam [4:0] OP5_OP_32 = 5'b01110;
               localparam [4:0] OP5_64B = 5'b01111;
               localparam [4:0] OP5_MADD = 5'b10000;
               localparam [4:0] OP5_MSUB = 5'b10001;
               localparam [4:0] OP5_NMSUB = 5'b10010;
               localparam [4:0] OP5_NMADD = 5'b10011;
               localparam [4:0] OP5_OP_FP = 5'b10100;  // (R-type, but rs2 = const for some, based on funct7 which doesn't exist for I-type?? R-type w/ ignored R2?)
               localparam [4:0] OP5_RESERVED_1 = 5'b10101;
               localparam [4:0] OP5_CUSTOM_2_RV128 = 5'b10110;
               localparam [4:0] OP5_48B2 = 5'b10111;
               localparam [4:0] OP5_BRANCH = 5'b11000;
               localparam [4:0] OP5_JALR = 5'b11001;
               localparam [4:0] OP5_RESERVED_2 = 5'b11010;
               localparam [4:0] OP5_JAL = 5'b11011;
               localparam [4:0] OP5_SYSTEM = 5'b11100;
               localparam [4:0] OP5_RESERVED_3 = 5'b11101;
               localparam [4:0] OP5_CUSTOM_3_RV128 = 5'b11110;
               localparam [4:0] OP5_80B = 5'b11111;
               
            /*SV_plus*/
               // Not sure these are ever used.
               localparam INSTR_TYPE_I_MASK = 0 | (1 << 5'b00000) | (1 << 5'b00001) | (1 << 5'b00100) | (1 << 5'b00110) | (1 << 5'b11001) | (1 << 5'b11100); localparam INSTR_TYPE_R_MASK = 0 | (1 << 5'b01100) | (1 << 5'b01110); localparam INSTR_TYPE_RI_MASK = 0 | (1 << 5'b01011) | (1 << 5'b10100); localparam INSTR_TYPE_R4_MASK = 0 | (1 << 5'b10000) | (1 << 5'b10001) | (1 << 5'b10010) | (1 << 5'b10011); localparam INSTR_TYPE_S_MASK = 0 | (1 << 5'b01000) | (1 << 5'b01001); localparam INSTR_TYPE_B_MASK = 0 | (1 << 5'b11000); localparam INSTR_TYPE_J_MASK = 0 | (1 << 5'b11011); localparam INSTR_TYPE_U_MASK = 0 | (1 << 5'b00101) | (1 << 5'b01101); localparam INSTR_TYPE___MASK = 0 | (1 << 5'b00010) | (1 << 5'b00011) | (1 << 5'b00111) | (1 << 5'b01010) | (1 << 5'b01111) | (1 << 5'b10101) | (1 << 5'b10110) | (1 << 5'b10111) | (1 << 5'b11010) | (1 << 5'b11101) | (1 << 5'b11110) | (1 << 5'b11111); 
               
            /*SV_plus*/
               // Instruction characterization.
               // (User ISA Manual 2.2, Table 19.2)
               // instr(type,  // (this is simply verified vs. op5)
               //       |  bit-width,
               //       |  |   extension, 
               //       |  |   |  opcode[6:2],  // (aka op5)
               //       |  |   |  |      func3,   // (if applicable)
               //       |  |   |  |      |    mnemonic)
               localparam [6:0] LUI_INSTR_OPCODE = 7'b0110111;
               localparam [6:0] AUIPC_INSTR_OPCODE = 7'b0010111;
               localparam [6:0] JAL_INSTR_OPCODE = 7'b1101111;
               localparam [6:0] JALR_INSTR_OPCODE = 7'b1100111; localparam [2:0] JALR_INSTR_FUNCT3 = 3'b000;
               localparam [6:0] BEQ_INSTR_OPCODE = 7'b1100011; localparam [2:0] BEQ_INSTR_FUNCT3 = 3'b000;
               localparam [6:0] BNE_INSTR_OPCODE = 7'b1100011; localparam [2:0] BNE_INSTR_FUNCT3 = 3'b001;
               localparam [6:0] BLT_INSTR_OPCODE = 7'b1100011; localparam [2:0] BLT_INSTR_FUNCT3 = 3'b100;
               localparam [6:0] BGE_INSTR_OPCODE = 7'b1100011; localparam [2:0] BGE_INSTR_FUNCT3 = 3'b101;
               localparam [6:0] BLTU_INSTR_OPCODE = 7'b1100011; localparam [2:0] BLTU_INSTR_FUNCT3 = 3'b110;
               localparam [6:0] BGEU_INSTR_OPCODE = 7'b1100011; localparam [2:0] BGEU_INSTR_FUNCT3 = 3'b111;
               localparam [6:0] LB_INSTR_OPCODE = 7'b0000011; localparam [2:0] LB_INSTR_FUNCT3 = 3'b000;
               localparam [6:0] LH_INSTR_OPCODE = 7'b0000011; localparam [2:0] LH_INSTR_FUNCT3 = 3'b001;
               localparam [6:0] LW_INSTR_OPCODE = 7'b0000011; localparam [2:0] LW_INSTR_FUNCT3 = 3'b010;
               localparam [6:0] LBU_INSTR_OPCODE = 7'b0000011; localparam [2:0] LBU_INSTR_FUNCT3 = 3'b100;
               localparam [6:0] LHU_INSTR_OPCODE = 7'b0000011; localparam [2:0] LHU_INSTR_FUNCT3 = 3'b101;
               localparam [6:0] SB_INSTR_OPCODE = 7'b0100011; localparam [2:0] SB_INSTR_FUNCT3 = 3'b000;
               localparam [6:0] SH_INSTR_OPCODE = 7'b0100011; localparam [2:0] SH_INSTR_FUNCT3 = 3'b001;
               localparam [6:0] SW_INSTR_OPCODE = 7'b0100011; localparam [2:0] SW_INSTR_FUNCT3 = 3'b010;
               localparam [6:0] ADDI_INSTR_OPCODE = 7'b0010011; localparam [2:0] ADDI_INSTR_FUNCT3 = 3'b000;
               localparam [6:0] SLTI_INSTR_OPCODE = 7'b0010011; localparam [2:0] SLTI_INSTR_FUNCT3 = 3'b010;
               localparam [6:0] SLTIU_INSTR_OPCODE = 7'b0010011; localparam [2:0] SLTIU_INSTR_FUNCT3 = 3'b011;
               localparam [6:0] XORI_INSTR_OPCODE = 7'b0010011; localparam [2:0] XORI_INSTR_FUNCT3 = 3'b100;
               localparam [6:0] ORI_INSTR_OPCODE = 7'b0010011; localparam [2:0] ORI_INSTR_FUNCT3 = 3'b110;
               localparam [6:0] ANDI_INSTR_OPCODE = 7'b0010011; localparam [2:0] ANDI_INSTR_FUNCT3 = 3'b111;
               localparam [6:0] SLLI_INSTR_OPCODE = 7'b0010011; localparam [2:0] SLLI_INSTR_FUNCT3 = 3'b001;
               localparam [6:0] SRLI_SRAI_INSTR_OPCODE = 7'b0010011; localparam [2:0] SRLI_SRAI_INSTR_FUNCT3 = 3'b101;  // Two instructions distinguished by an immediate bit, treated as a single instruction.
               localparam [6:0] ADD_SUB_INSTR_OPCODE = 7'b0110011; localparam [2:0] ADD_SUB_INSTR_FUNCT3 = 3'b000;  // Treated as a single instruction.
               localparam [6:0] SLL_INSTR_OPCODE = 7'b0110011; localparam [2:0] SLL_INSTR_FUNCT3 = 3'b001;
               localparam [6:0] SLT_INSTR_OPCODE = 7'b0110011; localparam [2:0] SLT_INSTR_FUNCT3 = 3'b010;
               localparam [6:0] SLTU_INSTR_OPCODE = 7'b0110011; localparam [2:0] SLTU_INSTR_FUNCT3 = 3'b011;
               localparam [6:0] XOR_INSTR_OPCODE = 7'b0110011; localparam [2:0] XOR_INSTR_FUNCT3 = 3'b100;
               localparam [6:0] SRL_SRA_INSTR_OPCODE = 7'b0110011; localparam [2:0] SRL_SRA_INSTR_FUNCT3 = 3'b101;  // Treated as a single instruction.
               localparam [6:0] OR_INSTR_OPCODE = 7'b0110011; localparam [2:0] OR_INSTR_FUNCT3 = 3'b110;
               localparam [6:0] AND_INSTR_OPCODE = 7'b0110011; localparam [2:0] AND_INSTR_FUNCT3 = 3'b111;
               //m4_instr(_, 32, I, 00011, 000, FENCE)
               //m4_instr(_, 32, I, 00011, 001, FENCE_I)
               //m4_instr(_, 32, I, 11100, 000, ECALL_EBREAK)  // Two instructions distinguished by an immediate bit, treated as a single instruction.
               localparam [6:0] CSRRW_INSTR_OPCODE = 7'b1110011; localparam [2:0] CSRRW_INSTR_FUNCT3 = 3'b001;
               localparam [6:0] CSRRS_INSTR_OPCODE = 7'b1110011; localparam [2:0] CSRRS_INSTR_FUNCT3 = 3'b010;
               localparam [6:0] CSRRC_INSTR_OPCODE = 7'b1110011; localparam [2:0] CSRRC_INSTR_FUNCT3 = 3'b011;
               localparam [6:0] CSRRWI_INSTR_OPCODE = 7'b1110011; localparam [2:0] CSRRWI_INSTR_FUNCT3 = 3'b101;
               localparam [6:0] CSRRSI_INSTR_OPCODE = 7'b1110011; localparam [2:0] CSRRSI_INSTR_FUNCT3 = 3'b110;
               localparam [6:0] CSRRCI_INSTR_OPCODE = 7'b1110011; localparam [2:0] CSRRCI_INSTR_FUNCT3 = 3'b111;
               
               
               
               
                 // Two instructions distinguished by an immediate bit, treated as a single instruction.
               
               
                 // Two instructions distinguished by an immediate bit, treated as a single instruction.
                 // Two instructions distinguished by an immediate bit, treated as a single instruction.
               
                 // Two instructions distinguished by an immediate bit, treated as a single instruction.
               
               
               
               
               
               
               
               
               
               
               
               
               
               // RV32A and RV64A
               // NOT IMPLEMENTED. These are distinct in the func7 field.
               // RV32F and RV64F
               // NOT IMPLEMENTED.
               // RV32D and RV64D
               // NOT IMPLEMENTED.
         
         
            // ^---------------------
            
         //_\end_source
   
      
      // The program in an instruction memory.
      /*SV_plus*/
         //logic [31:0] instrs [0:11-1];
      //_\source <builtin> 1   // Instantiated from warp-v_5-stage.tlv, 11 as: m4+indirect(M4_isa['_cnt10_prog'])
         //_\source ./warpv.tlv 1087   // Instantiated from built-in definition.
            
            /*SV_plus*/
               logic [40*8-1:0] instr_strs [0:11];
               
               // /=====================\
               // | Count to 10 Program |
               // \=====================/
               //
               
               // Add 1,2,3,...,10 (in that order).
               // Store incremental results in memory locations 0..9. (1, 3, 6, 10, ...)
               //
               // Regs:
               // 1: cnt
               // 2: ten
               // 3: out
               // 4: tmp
               // 5: offset
               // 6: store addr
               
/*               assign instrs = '{
                  {12'b0, 5'd0, ORI_INSTR_FUNCT3, 5'd6, ORI_INSTR_OPCODE},        //     store_addr = 0
                  {12'b1, 5'd0, ORI_INSTR_FUNCT3, 5'd1, ORI_INSTR_OPCODE},        //     cnt = 1
                  {12'b1010, 5'd0, ORI_INSTR_FUNCT3, 5'd2, ORI_INSTR_OPCODE},     //     ten = 10
                  {12'b0, 5'd0, ORI_INSTR_FUNCT3, 5'd3, ORI_INSTR_OPCODE},        //     out = 0
                  {7'b0, 5'd3, 5'd1, ADD_SUB_INSTR_FUNCT3, 5'd3, ADD_SUB_INSTR_OPCODE},       //  -> out += cnt
                  {7'b0000000, 5'd3, 5'd6, SW_INSTR_FUNCT3, 5'b00000, SW_INSTR_OPCODE},         //     store out at store_addr
                  {12'b1, 5'd1, ADDI_INSTR_FUNCT3, 5'd1, ADDI_INSTR_OPCODE},       //     cnt ++
                  {12'b100, 5'd6, ADDI_INSTR_FUNCT3, 5'd6, ADDI_INSTR_OPCODE},     //     store_addr++
                  {1'b1, 6'b111111, 5'd2, 5'd1, BLT_INSTR_FUNCT3, 4'b1000, 1'b1, BLT_INSTR_OPCODE}, //  ^- branch back if cnt < 10
                  {12'b111111111100, 5'd6, LW_INSTR_FUNCT3, 5'd4, LW_INSTR_OPCODE}, //     load the final value into tmp
                  {1'b1, 6'b111110, 5'd2, 5'd1, BGE_INSTR_FUNCT3, 4'b1010, 1'b1, BGE_INSTR_OPCODE}  //     TERMINATE by branching to -1
               };*/
               
               assign instr_strs = '{ "(I) ORI r6,r0,0                         ",  "(I) ORI r1,r0,1                         ",  "(I) ORI r2,r0,1010                      ",  "(I) ORI r3,r0,0                         ",  "(R) ADD_SUB r3,r1,r3                    ",  "(S) SW r6,r3,0                          ",  "(I) ADDI r1,r1,1                        ",  "(I) ADDI r6,r6,100                      ",  "(B) BLT r1,r2,1111111110000             ",  "(I) LW r4,r6,111111111100               ",  "(B) BGE r1,r2,1111111010100             ",  "END                                     "};
            //_|fetch
               for (instrs = 0; instrs <= 11; instrs++) begin : L1_FETCH_Instrs //_/instrs
                  //_@0  // whatever the fetch stage is.
                     assign FETCH_Instrs_instr_a0[instrs][31:0] =
                        (instrs == 0 ) ? {12'b0, 5'd0, ORI_INSTR_FUNCT3, 5'd6, ORI_INSTR_OPCODE} :
                        (instrs == 1 ) ? {12'b1, 5'd0, ORI_INSTR_FUNCT3, 5'd1, ORI_INSTR_OPCODE} :
                        (instrs == 2 ) ? {12'b1010, 5'd0, ORI_INSTR_FUNCT3, 5'd2, ORI_INSTR_OPCODE} :
                        (instrs == 3 ) ? {12'b0, 5'd0, ORI_INSTR_FUNCT3, 5'd3, ORI_INSTR_OPCODE} :
                        (instrs == 4 ) ? {7'b0, 5'd3, 5'd1, ADD_SUB_INSTR_FUNCT3, 5'd3, ADD_SUB_INSTR_OPCODE} :
                        (instrs == 5 ) ? {7'b0000000, 5'd3, 5'd6, SW_INSTR_FUNCT3, 5'b00000, SW_INSTR_OPCODE} :
                        (instrs == 6 ) ? {12'b1, 5'd1, ADDI_INSTR_FUNCT3, 5'd1, ADDI_INSTR_OPCODE} :
                        (instrs == 7 ) ? {12'b100, 5'd6, ADDI_INSTR_FUNCT3, 5'd6, ADDI_INSTR_OPCODE} :
                        (instrs == 8 ) ? {1'b1, 6'b111111, 5'd2, 5'd1, BLT_INSTR_FUNCT3, 4'b1000, 1'b1, BLT_INSTR_OPCODE} :
                        (instrs == 9 ) ? {12'b111111111100, 5'd6, LW_INSTR_FUNCT3, 5'd4, LW_INSTR_OPCODE} :
                        (instrs == 10 ) ?{1'b1, 6'b111110, 5'd2, 5'd1, BGE_INSTR_FUNCT3, 4'b1010, 1'b1, BGE_INSTR_OPCODE}: 32'b0;
                                       
               end
            
         //_\end_source
      
   
   
      // /=========\
      // | The CPU |
      // \=========/
   
      //_|fetch
         //_/instr
            // Provide a longer reset to cover the pipeline depth.
            //_@-1
               assign FETCH_Instr_Cnt_n2[7:0] = reset        ? 8'b0 :       // reset
                            FETCH_Instr_Cnt_n1 == 8'hFF ? 8'hFF :      // max out to avoid wrapping
                                            FETCH_Instr_Cnt_n1 + 8'b1; // increment
               assign FETCH_Instr_reset_n1 = reset || FETCH_Instr_Cnt_n1 < 5;
            
            //_@0
               assign FETCH_Instr_fetch_a0 = ! FETCH_Instr_reset_a0;  // always fetch
               //_?$fetch
   
                  // =====
                  // Fetch
                  // =====
   
                  // Fetch the raw instruction from program memory (or, for formal, tie it off).
                  
                  
                  
                  assign FETCH_Instr_raw_a0[31:0] = FETCH_Instrs_instr_a0[FETCH_Instr_Pc_a0[5:2]];
                  
            //_@0
               
               // ========
               // Overview
               // ========
               
               // Terminology:
               //
               // Instruction: An instruction, as viewed by the CPU pipeline (i.e. ld and returning_ld are separate instructions,
               //              and the returning_ld and the instruction it clobbers are one in the same).
               // ISA Instruction: An instruction, as defined by the ISA.
               // Good-Path (vs. Bad-Path): On the proper flow of execution of the program, excluding aborted instructions.
               // Path (of an instruction): The sequence of instructions that led to a particular instruction.
               // Current Path: The sequence of instructions fetched by next-PC logic that are not known to be bad-path.
               // Redirect: Adjust the PC from the predicted next-PC.
               // Redirect Shadow: Between the instruction causing the redirect and the redirect target instruction.
               // Bubbles: The cycles in the redirect shadow.
               // Commit: Results are made visible to subsequent instructions.
               // Abort: Do not commit. All aborts are also redirects and put the instruction on bad path. Non-aborting
               //        redirects do not mark the triggering instruction as bad-path. Aborts mask future redirects on the
               //        aborted instruction.
               // Retire: Commit results of an ISA instruction.
               
               // Control flow:
               //
               // Redirects include (earliest to latest):
               //   o Returning load: (aborting) A returning load clobbers an instruction and takes its slot, resulting in a
               //                     one-cycle redirect to repeat the clobbered instruction.
               //   o Predict-taken branch: A predicted-taken branch must determine the target before it can redirect the PC.
               //                           (This might be followed up by a mispredition.)
               //   o Replay: (aborting) Replay the same instruction (because a source register is pending (awaiting a returning_ld))
               //   o Jump: A jump instruction.
               //   o Mispredicted branch: A branch condition was mispredicted.
               //   o Aborting traps: (aborting) illegal instructions, others?
               //   o Non-aborting traps: misaligned PC target
               
               // ==============
               // Redirect Logic
               // ==============
                               
               // PC logic will redirect the PC for conditions on current-path instructions. PC logic keeps track of which
               // instructions are on the current path with a $GoodPathMask. $GoodPathMask[n] of an instruction indicates
               // whether the instruction n instructions prior to this instruction is on its path.
               //
               //                 $GoodPathMask for Redir'edX => {o,X,o,o,y,y,o,o} == {1,1,1,1,0,0,1,1}
               // Waterfall View: |
               //                 V
               // 0)       oooooooo                  Good-path
               // 1) InstX  ooooooXo  (Non-aborting) Good-path
               // 2)         ooooooxx
               // 3) InstY    ooYyyxxx  (Aborting)
               // 4) InstZ     ooyyxZxx
               // 5) Redir'edY  oyyxxxxx
               // 6) TargetY     ooxxxxxx
               // 7) Redir'edX    oxxxxxxx
               // 8) TargetX       oooooooo          Good-path
               // 9) Not redir'edZ  oooooooo         Good-path
               //
               // Above depicts a waterfall diagram where three triggering redirection conditions X, Y, and Z are detected on three different
               // instructions. A trigger in the 1st depicted stage, M4_NEXT_PC_STAGE, results in a zero-bubble redirect so it would be
               // a condition that is factored directly into the next-PC logic of the triggering instruction, and it would have
               // no impact on the $GoodPathMask.
               //
               // Waveform View:
               //
               //   Inst 0123456789
               //        ---------- /
               // GPM[7]        ooxxxxxxoo
               // GPM[6]       oXxxxxxxoo
               // GPM[5]      oooxZxxxoo
               // GPM[4]     oooyxxxxoo
               // GPM[3]    oooyyxxxoo
               // GPM[2]   oooYyyxxoo
               // GPM[1]  oooooyoxoo
               // GPM[0] oooooooooo
               //          /
               //         Triggers for Inst 3
               //
               // In the waveform view, the mask shifts up each cycle, as instructions age, and trigger conditions mask instructions
               // in the shadow, down to the redirect target (GPM[0]).
               //
               // Terminology:
               //   Triggering instruction: The instruction on which the condition is detected.
               //   Redirected instruction: The instruction whose next PC is redirected.
               //   Redirection target instruction: The first new-path instruction resulting from the redirection.
               //
               // Above, Y redirects first, though it is for a later instruction than X. The redirections for X and Y are taken
               // because their instructions are on the path of the redirected instructions. Z is not on the path of its
               // potentially-redirected instruction, so no redirection happens.
               //
               // For simultaneous conditions on different instructions, the PC must redirect to the earlier instruction's
               // redirect target, so later-stage redirects take priority in the PC-mux.
               //
               // Aborting redirects result in the aborting instruction being marked as bad-path. Aborted instructions will
               // not commit. Subsequent redirect conditions on aborting instructions are ignored. (For conditions within the
               // same stage, this is accomplished by the PC-mux prioritization.)
               
               
               // Macros are defined elsewhere based on the ordered set of conditions that generate code here.
               
               // Redirect Shadow
               // A mask of stages ahead of this one (older) in which instructions are on the path of this instruction.
               // Index 1 is ahead by 1, etc.
               // In the example above, $GoodPathMask for Redir'edX == {0,0,0,0,1,1,0,0}
               //     (Looking up in the waterfall diagram from its first "o", in reverse order {o,X,o,o,y,y,o,o}.)
               // The LSB is fetch-valid. It only exists for m4_valid_as_of macro.
               assign FETCH_Instr_next_good_path_mask_a0[1+1:0] =
                  // Shift up and mask w/ redirect conditions.
                  {FETCH_Instr_GoodPathMask_a0[1:0]
                   // & terms for each condition (order doesn't matter since masks are the same within a cycle)
                    & ((FETCH_Instr_returning_ld_a0 && !(1'b0) && FETCH_Instr_GoodPathMask_a0[0]) ? {{1{1'b1}}, {1{1'b0}}} : {2{1'b1}}) & ((FETCH_Instr_replay_a0 && !(1'b0 || FETCH_Instr_returning_ld_a0) && FETCH_Instr_GoodPathMask_a0[0]) ? {{1{1'b1}}, {1{1'b0}}} : {2{1'b1}}) & ((FETCH_Instr_jump_a0 && !(1'b0 || FETCH_Instr_returning_ld_a0 || FETCH_Instr_replay_a0) && FETCH_Instr_GoodPathMask_a0[0]) ? {{2{1'b1}}, {0{1'b0}}} : {2{1'b1}}) & ((FETCH_Instr_mispred_branch_a0 && !(1'b0 || FETCH_Instr_returning_ld_a0 || FETCH_Instr_replay_a0) && FETCH_Instr_GoodPathMask_a0[0]) ? {{2{1'b1}}, {0{1'b0}}} : {2{1'b1}}) & ((FETCH_Instr_indirect_jump_a0 && !(1'b0 || FETCH_Instr_returning_ld_a0 || FETCH_Instr_replay_a0) && FETCH_Instr_GoodPathMask_a0[0]) ? {{2{1'b1}}, {0{1'b0}}} : {2{1'b1}}) & ((FETCH_Instr_aborting_trap_a1 && !(1'b0 || FETCH_Instr_returning_ld_a1 || FETCH_Instr_replay_a1) && FETCH_Instr_GoodPathMask_a0[1]) ? {{0{1'b1}}, {2{1'b0}}} : {2{1'b1}}) & ((FETCH_Instr_non_aborting_trap_a1 && !(1'b0 || FETCH_Instr_returning_ld_a1 || FETCH_Instr_replay_a1 || FETCH_Instr_aborting_trap_a1) && FETCH_Instr_GoodPathMask_a0[1]) ? {{1{1'b1}}, {1{1'b0}}} : {2{1'b1}}),
                   1'b1}; // Shift in 1'b1 (fetch-valid).
               
               assign FETCH_Instr_GoodPathMask_n1[1+1:0] =
                  FETCH_Instr_reset_n1 ? 3'b0 :  // All bad-path (through self) on reset (next mask based on next reset).
                  FETCH_Instr_next_good_path_mask_a0;
               
               
               
               
               
                  
                   
                   
               
                  
                  
               
               
               
               // A returning load clobbers the instruction.
               // (Could do this with lower latency. Right now it goes through memory pipeline $ANY, and
               //  it is non-speculative. Both could easily be fixed.)
               assign FETCH_Instr_returning_ld_a0 = MEM_Data_valid_ld_a1 && 1'b1;
               // Recirculate returning load.
               //_?$returning_ld
                  // This scope holds the original load for a returning load.
                  //_/original_ld
                     assign {FETCH_Instr_OriginalLd_addr_a0[1:0], FETCH_Instr_OriginalLd_dest_reg_a0[4:0], FETCH_Instr_OriginalLd_ld_st_half_a0, FETCH_Instr_OriginalLd_ld_st_word_a0, FETCH_Instr_OriginalLd_ld_value_a0[31:0], FETCH_Instr_OriginalLd_raw_funct3_a0[2]} = {MEM_Data_addr_a1, MEM_Data_dest_reg_a1, MEM_Data_ld_st_half_a1, MEM_Data_ld_st_word_a1, MEM_Data_ld_value_a1, MEM_Data_raw_funct3_a1};
                     for (src = 1; src <= 2; src++) begin : L1_FETCH_Instr_OriginalLd_Src //_/src

                        // For $dummy.
                        logic L1_dummy_a0;

                        assign {L1_dummy_a0} = {L1_MEM_Data_Src[src].L1_dummy_a1};
                     end
               
               // Next PC
               assign FETCH_Instr_Pc_n1[31:2] =
                  FETCH_Instr_reset_a0 ? 30'b0 :
                  // ? : terms for each condition (order does matter)
                  (FETCH_Instr_non_aborting_trap_a1 && !(1'b0 || FETCH_Instr_returning_ld_a1 || FETCH_Instr_replay_a1 || FETCH_Instr_aborting_trap_a1) && FETCH_Instr_GoodPathMask_a0[1]) ? FETCH_Instr_trap_target_a1 : (FETCH_Instr_aborting_trap_a1 && !(1'b0 || FETCH_Instr_returning_ld_a1 || FETCH_Instr_replay_a1) && FETCH_Instr_GoodPathMask_a0[1]) ? FETCH_Instr_trap_target_a1 : (FETCH_Instr_indirect_jump_a0 && !(1'b0 || FETCH_Instr_returning_ld_a0 || FETCH_Instr_replay_a0) && FETCH_Instr_GoodPathMask_a0[0]) ? FETCH_Instr_indirect_jump_target_a0 : (FETCH_Instr_mispred_branch_a0 && !(1'b0 || FETCH_Instr_returning_ld_a0 || FETCH_Instr_replay_a0) && FETCH_Instr_GoodPathMask_a0[0]) ? FETCH_Instr_branch_redir_pc_a0 : (FETCH_Instr_jump_a0 && !(1'b0 || FETCH_Instr_returning_ld_a0 || FETCH_Instr_replay_a0) && FETCH_Instr_GoodPathMask_a0[0]) ? FETCH_Instr_jump_target_a0 : (FETCH_Instr_replay_a0 && !(1'b0 || FETCH_Instr_returning_ld_a0) && FETCH_Instr_GoodPathMask_a0[0]) ? FETCH_Instr_Pc_a0 : (FETCH_Instr_returning_ld_a0 && !(1'b0) && FETCH_Instr_GoodPathMask_a0[0]) ? FETCH_Instr_Pc_a0 :        
                           FETCH_Instr_Pc_a0 + 30'b1;
            
            //_@0
   
               // ======
               // DECODE
               // ======
   
               // Decode of the fetched instruction
               assign FETCH_Instr_valid_decode_a0 = FETCH_Instr_fetch_a0;  // Always decode if we fetch.
               assign FETCH_Instr_valid_decode_branch_a0 = FETCH_Instr_valid_decode_a0 && FETCH_Instr_branch_a0;
               //_\source <builtin> 1   // Instantiated from warp-v_5-stage.tlv, 1962 as: m4+indirect(M4_isa['_decode'])
                  //_\source ./warpv.tlv 1384   // Instantiated from built-in definition.
                     // TODO: ?$valid_<stage> conditioning should be replaced by use of m4_valid_as_of(M4_BLAH_STAGE).
                     //_?$valid_decode
                  
                        // =================================
                  
                        // Extract fields of $raw (instruction) into $raw_<field>[x:0].
                        assign {FETCH_Instr_raw_funct7_a0[6:0], FETCH_Instr_raw_rs2_a0[4:0], FETCH_Instr_raw_rs1_a0[4:0], FETCH_Instr_raw_funct3_a0[2:0], FETCH_Instr_raw_rd_a0[4:0], FETCH_Instr_raw_op5_a0[4:0], FETCH_Instr_raw_op2_a0[1:0]} = FETCH_Instr_raw_a0;
                        `BOGUS_USE(FETCH_Instr_raw_funct7_a0 FETCH_Instr_raw_op2_a0)  // Delete once its used.
                        // Extract immediate fields into type-specific signals.
                        // (User ISA Manual 2.2, Fig. 2.4)
                        assign FETCH_Instr_raw_i_imm_a0[31:0] = {{21{FETCH_Instr_raw_a0[31]}}, FETCH_Instr_raw_a0[30:20]};
                        assign FETCH_Instr_raw_s_imm_a0[31:0] = {{21{FETCH_Instr_raw_a0[31]}}, FETCH_Instr_raw_a0[30:25], FETCH_Instr_raw_a0[11:7]};
                        assign FETCH_Instr_raw_b_imm_a0[31:0] = {{20{FETCH_Instr_raw_a0[31]}}, FETCH_Instr_raw_a0[7], FETCH_Instr_raw_a0[30:25], FETCH_Instr_raw_a0[11:8], 1'b0};
                        assign FETCH_Instr_raw_u_imm_a0[31:0] = {FETCH_Instr_raw_a0[31:12], {12{1'b0}}};
                        assign FETCH_Instr_raw_j_imm_a0[31:0] = {{12{FETCH_Instr_raw_a0[31]}}, FETCH_Instr_raw_a0[19:12], FETCH_Instr_raw_a0[20], FETCH_Instr_raw_a0[30:21], 1'b0};
                        // Extract other type/instruction-specific fields.
                        assign FETCH_Instr_raw_shamt_a0[6:0] = FETCH_Instr_raw_a0[26:20];
                        assign FETCH_Instr_raw_aq_a0 = FETCH_Instr_raw_a0[26];
                        assign FETCH_Instr_raw_rl_a0 = FETCH_Instr_raw_a0[25];
                        assign FETCH_Instr_raw_rs3_a0[4:0] = FETCH_Instr_raw_a0[31:27];
                        assign FETCH_Instr_raw_rm_a0[2:0] = FETCH_Instr_raw_funct3_a0;
                        `BOGUS_USE(FETCH_Instr_raw_shamt_a0 FETCH_Instr_raw_aq_a0 FETCH_Instr_raw_rl_a0 FETCH_Instr_raw_rs3_a0 FETCH_Instr_raw_rm_a0)  // Avoid "unused" messages. Remove these as they become used.
                  
                        // Instruction type decode
                        /*SV_plus*/
                           assign FETCH_Instr_is_i_type_a0 = INSTR_TYPE_I_MASK[FETCH_Instr_raw_op5_a0]; assign FETCH_Instr_is_r_type_a0 = INSTR_TYPE_R_MASK[FETCH_Instr_raw_op5_a0]; assign FETCH_Instr_is_ri_type_a0 = INSTR_TYPE_RI_MASK[FETCH_Instr_raw_op5_a0]; assign FETCH_Instr_is_r4_type_a0 = INSTR_TYPE_R4_MASK[FETCH_Instr_raw_op5_a0]; assign FETCH_Instr_is_s_type_a0 = INSTR_TYPE_S_MASK[FETCH_Instr_raw_op5_a0]; assign FETCH_Instr_is_b_type_a0 = INSTR_TYPE_B_MASK[FETCH_Instr_raw_op5_a0]; assign FETCH_Instr_is_j_type_a0 = INSTR_TYPE_J_MASK[FETCH_Instr_raw_op5_a0]; assign FETCH_Instr_is_u_type_a0 = INSTR_TYPE_U_MASK[FETCH_Instr_raw_op5_a0]; assign FETCH_Instr_is___type_a0 = INSTR_TYPE___MASK[FETCH_Instr_raw_op5_a0]; 
                  
                        // Instruction decode.
                        //_\source ./warpv.tlv 1376   // Instantiated from warp-v_5-stage.tlv, 1413 as: m4+riscv_decode_expr()
                           assign FETCH_Instr_is_lui_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01101;
                           assign FETCH_Instr_is_auipc_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00101;
                           assign FETCH_Instr_is_jal_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11011;
                           assign FETCH_Instr_is_jalr_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11001 && FETCH_Instr_raw_funct3_a0 == 3'b000;
                           assign FETCH_Instr_is_beq_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11000 && FETCH_Instr_raw_funct3_a0 == 3'b000;
                           assign FETCH_Instr_is_bne_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11000 && FETCH_Instr_raw_funct3_a0 == 3'b001;
                           assign FETCH_Instr_is_blt_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11000 && FETCH_Instr_raw_funct3_a0 == 3'b100;
                           assign FETCH_Instr_is_bge_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11000 && FETCH_Instr_raw_funct3_a0 == 3'b101;
                           assign FETCH_Instr_is_bltu_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11000 && FETCH_Instr_raw_funct3_a0 == 3'b110;
                           assign FETCH_Instr_is_bgeu_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11000 && FETCH_Instr_raw_funct3_a0 == 3'b111;
                           assign FETCH_Instr_is_lb_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00000 && FETCH_Instr_raw_funct3_a0 == 3'b000;
                           assign FETCH_Instr_is_lh_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00000 && FETCH_Instr_raw_funct3_a0 == 3'b001;
                           assign FETCH_Instr_is_lw_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00000 && FETCH_Instr_raw_funct3_a0 == 3'b010;
                           assign FETCH_Instr_is_lbu_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00000 && FETCH_Instr_raw_funct3_a0 == 3'b100;
                           assign FETCH_Instr_is_lhu_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00000 && FETCH_Instr_raw_funct3_a0 == 3'b101;
                           assign FETCH_Instr_is_sb_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01000 && FETCH_Instr_raw_funct3_a0 == 3'b000;
                           assign FETCH_Instr_is_sh_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01000 && FETCH_Instr_raw_funct3_a0 == 3'b001;
                           assign FETCH_Instr_is_sw_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01000 && FETCH_Instr_raw_funct3_a0 == 3'b010;
                           assign FETCH_Instr_is_addi_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00100 && FETCH_Instr_raw_funct3_a0 == 3'b000;
                           assign FETCH_Instr_is_slti_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00100 && FETCH_Instr_raw_funct3_a0 == 3'b010;
                           assign FETCH_Instr_is_sltiu_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00100 && FETCH_Instr_raw_funct3_a0 == 3'b011;
                           assign FETCH_Instr_is_xori_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00100 && FETCH_Instr_raw_funct3_a0 == 3'b100;
                           assign FETCH_Instr_is_ori_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00100 && FETCH_Instr_raw_funct3_a0 == 3'b110;
                           assign FETCH_Instr_is_andi_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00100 && FETCH_Instr_raw_funct3_a0 == 3'b111;
                           assign FETCH_Instr_is_slli_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00100 && FETCH_Instr_raw_funct3_a0 == 3'b001;
                           assign FETCH_Instr_is_srli_srai_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b00100 && FETCH_Instr_raw_funct3_a0 == 3'b101;
                           assign FETCH_Instr_is_add_sub_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01100 && FETCH_Instr_raw_funct3_a0 == 3'b000;
                           assign FETCH_Instr_is_sll_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01100 && FETCH_Instr_raw_funct3_a0 == 3'b001;
                           assign FETCH_Instr_is_slt_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01100 && FETCH_Instr_raw_funct3_a0 == 3'b010;
                           assign FETCH_Instr_is_sltu_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01100 && FETCH_Instr_raw_funct3_a0 == 3'b011;
                           assign FETCH_Instr_is_xor_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01100 && FETCH_Instr_raw_funct3_a0 == 3'b100;
                           assign FETCH_Instr_is_srl_sra_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01100 && FETCH_Instr_raw_funct3_a0 == 3'b101;
                           assign FETCH_Instr_is_or_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01100 && FETCH_Instr_raw_funct3_a0 == 3'b110;
                           assign FETCH_Instr_is_and_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b01100 && FETCH_Instr_raw_funct3_a0 == 3'b111;
                           assign FETCH_Instr_is_csrrw_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11100 && FETCH_Instr_raw_funct3_a0 == 3'b001;
                           assign FETCH_Instr_is_csrrs_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11100 && FETCH_Instr_raw_funct3_a0 == 3'b010;
                           assign FETCH_Instr_is_csrrc_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11100 && FETCH_Instr_raw_funct3_a0 == 3'b011;
                           assign FETCH_Instr_is_csrrwi_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11100 && FETCH_Instr_raw_funct3_a0 == 3'b101;
                           assign FETCH_Instr_is_csrrsi_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11100 && FETCH_Instr_raw_funct3_a0 == 3'b110;
                           assign FETCH_Instr_is_csrrci_instr_a0 = FETCH_Instr_raw_op5_a0 == 5'b11100 && FETCH_Instr_raw_funct3_a0 == 3'b111;
                           
                        //_\end_source
                  
                        assign FETCH_Instr_illegal_a0 = 1'b1 && ! FETCH_Instr_is_lui_instr_a0 && ! FETCH_Instr_is_auipc_instr_a0 && ! FETCH_Instr_is_jal_instr_a0 && ! FETCH_Instr_is_jalr_instr_a0 && ! FETCH_Instr_is_beq_instr_a0 && ! FETCH_Instr_is_bne_instr_a0 && ! FETCH_Instr_is_blt_instr_a0 && ! FETCH_Instr_is_bge_instr_a0 && ! FETCH_Instr_is_bltu_instr_a0 && ! FETCH_Instr_is_bgeu_instr_a0 && ! FETCH_Instr_is_lb_instr_a0 && ! FETCH_Instr_is_lh_instr_a0 && ! FETCH_Instr_is_lw_instr_a0 && ! FETCH_Instr_is_lbu_instr_a0 && ! FETCH_Instr_is_lhu_instr_a0 && ! FETCH_Instr_is_sb_instr_a0 && ! FETCH_Instr_is_sh_instr_a0 && ! FETCH_Instr_is_sw_instr_a0 && ! FETCH_Instr_is_addi_instr_a0 && ! FETCH_Instr_is_slti_instr_a0 && ! FETCH_Instr_is_sltiu_instr_a0 && ! FETCH_Instr_is_xori_instr_a0 && ! FETCH_Instr_is_ori_instr_a0 && ! FETCH_Instr_is_andi_instr_a0 && ! FETCH_Instr_is_slli_instr_a0 && ! FETCH_Instr_is_srli_srai_instr_a0 && ! FETCH_Instr_is_add_sub_instr_a0 && ! FETCH_Instr_is_sll_instr_a0 && ! FETCH_Instr_is_slt_instr_a0 && ! FETCH_Instr_is_sltu_instr_a0 && ! FETCH_Instr_is_xor_instr_a0 && ! FETCH_Instr_is_srl_sra_instr_a0 && ! FETCH_Instr_is_or_instr_a0 && ! FETCH_Instr_is_and_instr_a0 && ! FETCH_Instr_is_csrrw_instr_a0 && ! FETCH_Instr_is_csrrs_instr_a0 && ! FETCH_Instr_is_csrrc_instr_a0 && ! FETCH_Instr_is_csrrwi_instr_a0 && ! FETCH_Instr_is_csrrsi_instr_a0 && ! FETCH_Instr_is_csrrci_instr_a0;
                        assign FETCH_Instr_conditional_branch_a0 = FETCH_Instr_is_b_type_a0;
                     assign FETCH_Instr_jump_a0 = FETCH_Instr_is_jal_instr_a0;  // "Jump" in RISC-V means unconditional. (JALR is a separate redirect condition.)
                     assign FETCH_Instr_branch_a0 = FETCH_Instr_is_b_type_a0;
                     assign FETCH_Instr_indirect_jump_a0 = FETCH_Instr_is_jalr_instr_a0;
                     //_?$valid_decode
                        assign FETCH_Instr_ld_a0 = FETCH_Instr_raw_a0[6:3] == 4'b0;
                        assign FETCH_Instr_st_a0 = FETCH_Instr_is_s_type_a0;
                        assign FETCH_Instr_ld_st_a0 = FETCH_Instr_ld_a0 || FETCH_Instr_st_a0;
                        assign FETCH_Instr_ld_st_word_a0 = FETCH_Instr_ld_st_a0 && (FETCH_Instr_raw_funct3_a0[1] == 1'b1);
                        assign FETCH_Instr_ld_st_half_a0 = FETCH_Instr_ld_st_a0 && (FETCH_Instr_raw_funct3_a0[1:0] == 2'b01);
                        //$ld_st_byte = $ld_st && ($raw_funct3[1:0] == 2'b00);
                        `BOGUS_USE(FETCH_Instr_is___type_a0 FETCH_Instr_is_u_type_a0)
                  
                        // Output signals.
                        for (src = 1; src <= 2; src++) begin : L1_FETCH_Instr_Src //_/src

                           // For $is_reg.
                           logic L1_is_reg_a0;

                           // For $reg.
                           logic [4:0] L1_reg_a0;

                           // Reg valid for this source, based on instruction type.
                           assign L1_is_reg_a0 = FETCH_Instr_is_r_type_a0 || FETCH_Instr_is_r4_type_a0 || (FETCH_Instr_is_i_type_a0 && (src == 1)) || FETCH_Instr_is_ri_type_a0 || FETCH_Instr_is_s_type_a0 || FETCH_Instr_is_b_type_a0;
                           assign L1_reg_a0[4:0] = (src == 1) ? FETCH_Instr_raw_rs1_a0 : FETCH_Instr_raw_rs2_a0;
                             
                        end
                        // For debug.
                        assign FETCH_Instr_mnemonic_a0[10*8-1:0] = FETCH_Instr_is_lui_instr_a0 ? "LUI       " : FETCH_Instr_is_auipc_instr_a0 ? "AUIPC     " : FETCH_Instr_is_jal_instr_a0 ? "JAL       " : FETCH_Instr_is_jalr_instr_a0 ? "JALR      " : FETCH_Instr_is_beq_instr_a0 ? "BEQ       " : FETCH_Instr_is_bne_instr_a0 ? "BNE       " : FETCH_Instr_is_blt_instr_a0 ? "BLT       " : FETCH_Instr_is_bge_instr_a0 ? "BGE       " : FETCH_Instr_is_bltu_instr_a0 ? "BLTU      " : FETCH_Instr_is_bgeu_instr_a0 ? "BGEU      " : FETCH_Instr_is_lb_instr_a0 ? "LB        " : FETCH_Instr_is_lh_instr_a0 ? "LH        " : FETCH_Instr_is_lw_instr_a0 ? "LW        " : FETCH_Instr_is_lbu_instr_a0 ? "LBU       " : FETCH_Instr_is_lhu_instr_a0 ? "LHU       " : FETCH_Instr_is_sb_instr_a0 ? "SB        " : FETCH_Instr_is_sh_instr_a0 ? "SH        " : FETCH_Instr_is_sw_instr_a0 ? "SW        " : FETCH_Instr_is_addi_instr_a0 ? "ADDI      " : FETCH_Instr_is_slti_instr_a0 ? "SLTI      " : FETCH_Instr_is_sltiu_instr_a0 ? "SLTIU     " : FETCH_Instr_is_xori_instr_a0 ? "XORI      " : FETCH_Instr_is_ori_instr_a0 ? "ORI       " : FETCH_Instr_is_andi_instr_a0 ? "ANDI      " : FETCH_Instr_is_slli_instr_a0 ? "SLLI      " : FETCH_Instr_is_srli_srai_instr_a0 ? "SRLI_SRAI " : FETCH_Instr_is_add_sub_instr_a0 ? "ADD_SUB   " : FETCH_Instr_is_sll_instr_a0 ? "SLL       " : FETCH_Instr_is_slt_instr_a0 ? "SLT       " : FETCH_Instr_is_sltu_instr_a0 ? "SLTU      " : FETCH_Instr_is_xor_instr_a0 ? "XOR       " : FETCH_Instr_is_srl_sra_instr_a0 ? "SRL_SRA   " : FETCH_Instr_is_or_instr_a0 ? "OR        " : FETCH_Instr_is_and_instr_a0 ? "AND       " : FETCH_Instr_is_csrrw_instr_a0 ? "CSRRW     " : FETCH_Instr_is_csrrs_instr_a0 ? "CSRRS     " : FETCH_Instr_is_csrrc_instr_a0 ? "CSRRC     " : FETCH_Instr_is_csrrwi_instr_a0 ? "CSRRWI    " : FETCH_Instr_is_csrrsi_instr_a0 ? "CSRRSI    " : FETCH_Instr_is_csrrci_instr_a0 ? "CSRRCI    " :  "ILLEGAL   ";
                        `BOGUS_USE(FETCH_Instr_mnemonic_a0)
                     // Condition signals must not themselves be conditioned (currently).
                     assign FETCH_Instr_dest_reg_a0[4:0] = FETCH_Instr_returning_ld_a0 ? FETCH_Instr_OriginalLd_dest_reg_a0 : FETCH_Instr_raw_rd_a0;
                     assign FETCH_Instr_dest_reg_valid_a0 = ((FETCH_Instr_valid_decode_a0 && ! FETCH_Instr_is_s_type_a0 && ! FETCH_Instr_is_b_type_a0) || FETCH_Instr_returning_ld_a0) &&
                                       | FETCH_Instr_dest_reg_a0;   // r0 not valid.
                     // Actually load.
                     assign FETCH_Instr_spec_ld_a0 = FETCH_Instr_valid_decode_a0 && FETCH_Instr_ld_a0;
                     
                  //_\end_source
            //_\source <builtin> 1   // Instantiated from warp-v_5-stage.tlv, 1963 as: m4+indirect(['branch_pred_']M4_BRANCH_PRED)
               //_\source ./warpv.tlv 1738   // Instantiated from built-in definition.
                  //_@0
                     assign FETCH_Instr_pred_taken_a0 = 1'b0;
               //_\end_source
            
            //_@0
               // Pending value to write to dest reg. Loads (not replaced by returning ld) write pending.
               assign FETCH_Instr_reg_wr_pending_a0 = FETCH_Instr_ld_a0 && ! FETCH_Instr_returning_ld_a0 && 1'b1;
               `BOGUS_USE(FETCH_Instr_reg_wr_pending_a0)  // Not used if no bypass and no pending.
               
               // ======
               // Reg Rd
               // ======
               
               // Obtain source register values and pending bit for source registers. Bypass up to 3
               // stages.
               // It is not necessary to bypass pending, as we could delay the replay, but we implement
               // bypass for performance.
               // Pending has an additional read for the dest register as we need to replay for write-after-write
               // hazard as well as write-after-read. To replay for dest write with the same timing, we must also
               // bypass the dest reg's pending bit.
               //_/regs
               for (src = 1; src <= 2; src++) begin : L1b_FETCH_Instr_Src //_/src

                  // For $dummy.
                  logic L1_dummy_a0;

                  // For $is_reg_condition.
                  logic L1_is_reg_condition_a0;

                  // For $pending.
                  logic L1_pending_a0;

                  // For $reg_value.
                  logic [31:0] L1_reg_value_a0;

                  assign L1_is_reg_condition_a0 = L1_FETCH_Instr_Src[src].L1_is_reg_a0 && FETCH_Instr_valid_decode_a0;  // Note: $is_reg can be set for RISC-V sr0.
                  //_?$is_reg_condition
                     assign {L1_reg_value_a0[31:0], L1_pending_a0} =
                        (L1_FETCH_Instr_Src[src].L1_reg_a0 == 5'b0) ? {32'b0, 1'b0} :  // Read r0 as 0 (not pending).
                        // Bypass stages. Both register and pending are bypassed.
                        // Bypassed registers must be from instructions that are good-path as of this instruction or are returning_ld.
                        
                        
                        
                        {FETCH_Instr_Regs_value_a0[L1_FETCH_Instr_Src[src].L1_reg_a0], FETCH_Instr_Regs_pending_a0[L1_FETCH_Instr_Src[src].L1_reg_a0]};
                  // Replay if this source register is pending.
                  assign FETCH_Instr_Src_replay_a0[src] = L1_is_reg_condition_a0 && L1_pending_a0;
                  assign L1_dummy_a0 = 1'b0;  // Dummy signal to pull through $ANY expressions when not building verification harness (since SandPiper currently complains about empty $ANY).
               end
               // Also replay for pending dest reg to keep writes in order. Bypass dest reg pending to support this.
               assign FETCH_Instr_is_dest_condition_a0 = FETCH_Instr_dest_reg_valid_a0 && FETCH_Instr_valid_decode_a0;  // Note, $dest_reg_valid is 0 for RISC-V sr0.
               //_?$is_dest_condition
                  assign FETCH_Instr_dest_pending_a0 =
                     (FETCH_Instr_dest_reg_a0 == 5'b0) ? 1'b0 :  // Read r0 as 0 (not pending). Not actually necessary, but it cuts off read of non-existent rs0, which might be an issue for formal verif tools.
                     // Bypass stages. Both register and pending are bypassed.
                     
                     
                     
                     FETCH_Instr_Regs_pending_a0[FETCH_Instr_dest_reg_a0];
               // Combine replay conditions for pending source or dest registers.
               assign FETCH_Instr_replay_a0 = | FETCH_Instr_Src_replay_a0 || (FETCH_Instr_is_dest_condition_a0 && FETCH_Instr_dest_pending_a0);
            
            
            // =======
            // Execute
            // =======
            //_\source <builtin> 1   // Instantiated from warp-v_5-stage.tlv, 2013 as: m4+indirect(M4_isa['_exe'], @M4_EXECUTE_STAGE, @M4_RESULT_STAGE)
               //_\source ./warpv.tlv 1445   // Instantiated from built-in definition.
                  //_@0
                     //_?$valid_decode_branch
                        assign FETCH_Instr_branch_target_a0[31:2] = FETCH_Instr_Pc_a0[31:2] + FETCH_Instr_raw_b_imm_a0[31:2];
                        assign FETCH_Instr_misaligned_pc_a0 = | FETCH_Instr_raw_b_imm_a0[1:0];
                     //_?$jump  // (JAL, not JALR)
                        assign FETCH_Instr_jump_target_a0[31:2] = FETCH_Instr_Pc_a0[31:2] + FETCH_Instr_raw_j_imm_a0[31:2];
                        assign FETCH_Instr_misaligned_jump_target_a0 = FETCH_Instr_raw_j_imm_a0[1];
                  //_@0
                     // Execution.
                     assign FETCH_Instr_valid_exe_a0 = FETCH_Instr_valid_decode_a0; // Execute if we decoded.
                     
                     // Compute results for each instruction, independent of decode (power-hungry, but fast).
                     //_?$valid_exe
                        assign FETCH_Instr_equal_a0 = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 == L1b_FETCH_Instr_Src[2].L1_reg_value_a0;
                     //_?$branch
                        assign FETCH_Instr_taken_a0 =
                           FETCH_Instr_is_j_type_a0 ||
                           (FETCH_Instr_is_beq_instr_a0 && FETCH_Instr_equal_a0) ||
                           (FETCH_Instr_is_bne_instr_a0 && ! FETCH_Instr_equal_a0) ||
                           ((FETCH_Instr_is_blt_instr_a0 || FETCH_Instr_is_bltu_instr_a0 || FETCH_Instr_is_bge_instr_a0 || FETCH_Instr_is_bgeu_instr_a0) &&
                            ((FETCH_Instr_is_bge_instr_a0 || FETCH_Instr_is_bgeu_instr_a0) ^
                             (({(FETCH_Instr_is_blt_instr_a0 ^ L1b_FETCH_Instr_Src[1].L1_reg_value_a0[31]), L1b_FETCH_Instr_Src[1].L1_reg_value_a0[31-1:0]} <
                              {(FETCH_Instr_is_blt_instr_a0 ^ L1b_FETCH_Instr_Src[2].L1_reg_value_a0[31]), L1b_FETCH_Instr_Src[2].L1_reg_value_a0[31-1:0]}) ^ ((L1b_FETCH_Instr_Src[1].L1_reg_value_a0[31] != L1b_FETCH_Instr_Src[2].L1_reg_value_a0[31]) & FETCH_Instr_is_bge_instr_a0)
                             )
                            )
                           );
                     //_?$indirect_jump  // (JALR)
                        assign FETCH_Instr_indirect_jump_full_target_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 + FETCH_Instr_raw_i_imm_a0;
                        assign FETCH_Instr_indirect_jump_target_a0[31:2] = FETCH_Instr_indirect_jump_full_target_a0[31:2];
                        assign FETCH_Instr_misaligned_indirect_jump_target_a0 = FETCH_Instr_indirect_jump_full_target_a0[1];
                     //_?$valid_exe
                        // Compute each individual instruction result, combined per-instruction by a macro.
                        
                        assign FETCH_Instr_lui_rslt_a0[31:0] = {FETCH_Instr_raw_u_imm_a0[31:12], 12'b0};
                        assign FETCH_Instr_auipc_rslt_a0[31:0] = {FETCH_Instr_Pc_a0, 2'b0} + FETCH_Instr_raw_u_imm_a0;
                        assign FETCH_Instr_jal_rslt_a0[31:0] = {FETCH_Instr_Pc_a0, 2'b0} + 4;
                        assign FETCH_Instr_jalr_rslt_a0[31:0] = {FETCH_Instr_Pc_a0, 2'b0} + 4;
                        // Load instructions. If returning ld is enabled, load instructions write no meaningful result, so we use zeros.
                        
                        assign FETCH_Instr_lb_rslt_a0[31:0] = 32'b0;
                        assign FETCH_Instr_lh_rslt_a0[31:0] = 32'b0;
                        assign FETCH_Instr_lw_rslt_a0[31:0] = 32'b0;
                        assign FETCH_Instr_lbu_rslt_a0[31:0] = 32'b0;
                        assign FETCH_Instr_lhu_rslt_a0[31:0] = 32'b0;
                        
                        
                        
                        
                        
                        
                        
                        assign FETCH_Instr_addi_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 + FETCH_Instr_raw_i_imm_a0;  // Note: this has its own adder; could share w/ add/sub.
                        assign FETCH_Instr_xori_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 ^ FETCH_Instr_raw_i_imm_a0;
                        assign FETCH_Instr_ori_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 | FETCH_Instr_raw_i_imm_a0;
                        assign FETCH_Instr_andi_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 & FETCH_Instr_raw_i_imm_a0;
                        assign FETCH_Instr_slli_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 << FETCH_Instr_raw_i_imm_a0[5:0];
                        assign FETCH_Instr_srli_intermediate_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 >> FETCH_Instr_raw_i_imm_a0[5:0];
                        assign FETCH_Instr_srai_intermediate_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0[31] ? FETCH_Instr_srli_intermediate_rslt_a0 | ((32'b0 - 1) << (32 - FETCH_Instr_raw_i_imm_a0[5:0]) ): FETCH_Instr_srli_intermediate_rslt_a0;
                        assign FETCH_Instr_sra_intermediate_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0[31] ? FETCH_Instr_srl_intermediate_rslt_a0 | ((32'b0 - 1) << (32 - L1b_FETCH_Instr_Src[2].L1_reg_value_a0[4:0]) ): FETCH_Instr_srl_intermediate_rslt_a0;
                        assign FETCH_Instr_srl_intermediate_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 >> L1b_FETCH_Instr_Src[2].L1_reg_value_a0[4:0];
                        assign FETCH_Instr_slti_rslt_a0[31:0] =  (L1b_FETCH_Instr_Src[1].L1_reg_value_a0[31] == FETCH_Instr_raw_i_imm_a0[31]) ? FETCH_Instr_sltiu_rslt_a0 : {31'b0,L1b_FETCH_Instr_Src[1].L1_reg_value_a0[31]};
                        assign FETCH_Instr_sltiu_rslt_a0[31:0] = (L1b_FETCH_Instr_Src[1].L1_reg_value_a0 < FETCH_Instr_raw_i_imm_a0) ? 1 : 0;
                        assign FETCH_Instr_srli_srai_rslt_a0[31:0] = (FETCH_Instr_raw_i_imm_a0[10] == 1) ? FETCH_Instr_srai_intermediate_rslt_a0 : FETCH_Instr_srli_intermediate_rslt_a0;
                        assign FETCH_Instr_add_sub_rslt_a0[31:0] =  (FETCH_Instr_raw_funct7_a0[5] == 1) ?  L1b_FETCH_Instr_Src[1].L1_reg_value_a0 - L1b_FETCH_Instr_Src[2].L1_reg_value_a0 : L1b_FETCH_Instr_Src[1].L1_reg_value_a0 + L1b_FETCH_Instr_Src[2].L1_reg_value_a0;
                        assign FETCH_Instr_sll_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 << L1b_FETCH_Instr_Src[2].L1_reg_value_a0[4:0];
                        assign FETCH_Instr_slt_rslt_a0[31:0] = (L1b_FETCH_Instr_Src[1].L1_reg_value_a0[31] == L1b_FETCH_Instr_Src[2].L1_reg_value_a0[31]) ? FETCH_Instr_sltu_rslt_a0 : {31'b0,L1b_FETCH_Instr_Src[1].L1_reg_value_a0[31]};
                        assign FETCH_Instr_sltu_rslt_a0[31:0] = (L1b_FETCH_Instr_Src[1].L1_reg_value_a0 < L1b_FETCH_Instr_Src[2].L1_reg_value_a0) ? 1 : 0;
                        assign FETCH_Instr_xor_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 ^ L1b_FETCH_Instr_Src[2].L1_reg_value_a0;
                        assign FETCH_Instr_srl_sra_rslt_a0[31:0] = (FETCH_Instr_raw_funct7_a0[5] == 1) ? FETCH_Instr_sra_intermediate_rslt_a0 : FETCH_Instr_srl_intermediate_rslt_a0;
                        assign FETCH_Instr_or_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 | L1b_FETCH_Instr_Src[2].L1_reg_value_a0;
                        assign FETCH_Instr_and_rslt_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 & L1b_FETCH_Instr_Src[2].L1_reg_value_a0;
                        // TODO: CSR read instructions have the same result expression. Synthesis might not optimize optimally.
                        assign FETCH_Instr_csrrw_rslt_a0[31:0]  = FETCH_Instr_is_csr_instreth_a0 ? FETCH_Instr_csr_instreth_a0 : FETCH_Instr_is_csr_instret_a0 ? FETCH_Instr_csr_instret_a0 : FETCH_Instr_is_csr_timeh_a0 ? FETCH_Instr_csr_timeh_a0 : FETCH_Instr_is_csr_time_a0 ? FETCH_Instr_csr_time_a0 : FETCH_Instr_is_csr_cycleh_a0 ? FETCH_Instr_csr_cycleh_a0 : FETCH_Instr_is_csr_cycle_a0 ? FETCH_Instr_csr_cycle_a0 : 32'bx;
                        assign FETCH_Instr_csrrs_rslt_a0[31:0]  = FETCH_Instr_is_csr_instreth_a0 ? FETCH_Instr_csr_instreth_a0 : FETCH_Instr_is_csr_instret_a0 ? FETCH_Instr_csr_instret_a0 : FETCH_Instr_is_csr_timeh_a0 ? FETCH_Instr_csr_timeh_a0 : FETCH_Instr_is_csr_time_a0 ? FETCH_Instr_csr_time_a0 : FETCH_Instr_is_csr_cycleh_a0 ? FETCH_Instr_csr_cycleh_a0 : FETCH_Instr_is_csr_cycle_a0 ? FETCH_Instr_csr_cycle_a0 : 32'bx;
                        assign FETCH_Instr_csrrc_rslt_a0[31:0]  = FETCH_Instr_is_csr_instreth_a0 ? FETCH_Instr_csr_instreth_a0 : FETCH_Instr_is_csr_instret_a0 ? FETCH_Instr_csr_instret_a0 : FETCH_Instr_is_csr_timeh_a0 ? FETCH_Instr_csr_timeh_a0 : FETCH_Instr_is_csr_time_a0 ? FETCH_Instr_csr_time_a0 : FETCH_Instr_is_csr_cycleh_a0 ? FETCH_Instr_csr_cycleh_a0 : FETCH_Instr_is_csr_cycle_a0 ? FETCH_Instr_csr_cycle_a0 : 32'bx;
                        assign FETCH_Instr_csrrwi_rslt_a0[31:0] = FETCH_Instr_is_csr_instreth_a0 ? FETCH_Instr_csr_instreth_a0 : FETCH_Instr_is_csr_instret_a0 ? FETCH_Instr_csr_instret_a0 : FETCH_Instr_is_csr_timeh_a0 ? FETCH_Instr_csr_timeh_a0 : FETCH_Instr_is_csr_time_a0 ? FETCH_Instr_csr_time_a0 : FETCH_Instr_is_csr_cycleh_a0 ? FETCH_Instr_csr_cycleh_a0 : FETCH_Instr_is_csr_cycle_a0 ? FETCH_Instr_csr_cycle_a0 : 32'bx;
                        assign FETCH_Instr_csrrsi_rslt_a0[31:0] = FETCH_Instr_is_csr_instreth_a0 ? FETCH_Instr_csr_instreth_a0 : FETCH_Instr_is_csr_instret_a0 ? FETCH_Instr_csr_instret_a0 : FETCH_Instr_is_csr_timeh_a0 ? FETCH_Instr_csr_timeh_a0 : FETCH_Instr_is_csr_time_a0 ? FETCH_Instr_csr_time_a0 : FETCH_Instr_is_csr_cycleh_a0 ? FETCH_Instr_csr_cycleh_a0 : FETCH_Instr_is_csr_cycle_a0 ? FETCH_Instr_csr_cycle_a0 : 32'bx;
                        assign FETCH_Instr_csrrci_rslt_a0[31:0] = FETCH_Instr_is_csr_instreth_a0 ? FETCH_Instr_csr_instreth_a0 : FETCH_Instr_is_csr_instret_a0 ? FETCH_Instr_csr_instret_a0 : FETCH_Instr_is_csr_timeh_a0 ? FETCH_Instr_csr_timeh_a0 : FETCH_Instr_is_csr_time_a0 ? FETCH_Instr_csr_time_a0 : FETCH_Instr_is_csr_cycleh_a0 ? FETCH_Instr_csr_cycleh_a0 : FETCH_Instr_is_csr_cycle_a0 ? FETCH_Instr_csr_cycle_a0 : 32'bx;
                        
                  // CSR logic
                  // ---------
                  //_\source ./warpv.tlv 1312   // Instantiated from warp-v_5-stage.tlv, 1527 as: m4+riscv_csrs((m4_csrs))
                     
                     //_\source ./warpv.tlv 1282   // Instantiated from warp-v_5-stage.tlv, 11 as: m4+riscv_csr(m4_echo(['m4_csr_']csr['_args']))
                        //--------------
                        // CSR CYCLE
                        //--------------
                        //_@0
                           assign FETCH_Instr_is_csr_cycle_a0 = FETCH_Instr_raw_a0[31:20] == 12'hC00;
                        //_@0
                           // CSR update. Counting on synthesis to optimize each bit, based on 32'b1.
                           
                           
                           // hw_wr_mask conditioned by hw_wr.
                           assign FETCH_Instr_csr_cycle_hw_wr_en_mask_a0[31:0] = {32{FETCH_Instr_csr_cycle_hw_wr_a0}} & FETCH_Instr_csr_cycle_hw_wr_mask_a0;
                           // The CSR value, updated by side-effect writes (if 1).
                           assign FETCH_Instr_upd_csr_cycle_a0[31:0] =
                                (FETCH_Instr_csr_cycle_hw_wr_en_mask_a0 & FETCH_Instr_csr_cycle_hw_wr_value_a0) | (! FETCH_Instr_csr_cycle_hw_wr_en_mask_a0 & FETCH_Instr_csr_cycle_a0);
                           // Next value of the CSR.
                           assign FETCH_Instr_csr_cycle_masked_wr_value_a0[31:0] =
                                FETCH_Instr_masked_csr_wr_value_a0[31:0] & 32'b1;
                           assign FETCH_Instr_csr_cycle_n1[31:0] =
                                FETCH_Instr_reset_a0 ? 32'b0 :
                                ((FETCH_Instr_is_csrrw_instr_a0 || FETCH_Instr_is_csrrwi_instr_a0) && FETCH_Instr_is_csr_cycle_a0)
                                       ? FETCH_Instr_csr_cycle_masked_wr_value_a0 | (FETCH_Instr_upd_csr_cycle_a0 & ! 32'b1) :
                                ((FETCH_Instr_is_csrrs_instr_a0 || FETCH_Instr_is_csrrsi_instr_a0) && FETCH_Instr_is_csr_cycle_a0)
                                       ? FETCH_Instr_upd_csr_cycle_a0 |   FETCH_Instr_csr_cycle_masked_wr_value_a0 :
                                ((FETCH_Instr_is_csrrc_instr_a0 || FETCH_Instr_is_csrrci_instr_a0) && FETCH_Instr_is_csr_cycle_a0)
                                       ? FETCH_Instr_upd_csr_cycle_a0 & ~ FETCH_Instr_csr_cycle_masked_wr_value_a0 :
                                // retain
                                         FETCH_Instr_upd_csr_cycle_a0;
                     //_\end_source
                     
                     //_\source ./warpv.tlv 1282   // Instantiated from warp-v_5-stage.tlv, 11 as: m4+riscv_csr(m4_echo(['m4_csr_']csr['_args']))
                        //--------------
                        // CSR CYCLEH
                        //--------------
                        //_@0
                           assign FETCH_Instr_is_csr_cycleh_a0 = FETCH_Instr_raw_a0[31:20] == 12'hC80;
                        //_@0
                           // CSR update. Counting on synthesis to optimize each bit, based on 32'b1.
                           
                           
                           // hw_wr_mask conditioned by hw_wr.
                           assign FETCH_Instr_csr_cycleh_hw_wr_en_mask_a0[31:0] = {32{FETCH_Instr_csr_cycleh_hw_wr_a0}} & FETCH_Instr_csr_cycleh_hw_wr_mask_a0;
                           // The CSR value, updated by side-effect writes (if 1).
                           assign FETCH_Instr_upd_csr_cycleh_a0[31:0] =
                                (FETCH_Instr_csr_cycleh_hw_wr_en_mask_a0 & FETCH_Instr_csr_cycleh_hw_wr_value_a0) | (! FETCH_Instr_csr_cycleh_hw_wr_en_mask_a0 & FETCH_Instr_csr_cycleh_a0);
                           // Next value of the CSR.
                           assign FETCH_Instr_csr_cycleh_masked_wr_value_a0[31:0] =
                                FETCH_Instr_masked_csr_wr_value_a0[31:0] & 32'b1;
                           assign FETCH_Instr_csr_cycleh_n1[31:0] =
                                FETCH_Instr_reset_a0 ? 32'b0 :
                                ((FETCH_Instr_is_csrrw_instr_a0 || FETCH_Instr_is_csrrwi_instr_a0) && FETCH_Instr_is_csr_cycleh_a0)
                                       ? FETCH_Instr_csr_cycleh_masked_wr_value_a0 | (FETCH_Instr_upd_csr_cycleh_a0 & ! 32'b1) :
                                ((FETCH_Instr_is_csrrs_instr_a0 || FETCH_Instr_is_csrrsi_instr_a0) && FETCH_Instr_is_csr_cycleh_a0)
                                       ? FETCH_Instr_upd_csr_cycleh_a0 |   FETCH_Instr_csr_cycleh_masked_wr_value_a0 :
                                ((FETCH_Instr_is_csrrc_instr_a0 || FETCH_Instr_is_csrrci_instr_a0) && FETCH_Instr_is_csr_cycleh_a0)
                                       ? FETCH_Instr_upd_csr_cycleh_a0 & ~ FETCH_Instr_csr_cycleh_masked_wr_value_a0 :
                                // retain
                                         FETCH_Instr_upd_csr_cycleh_a0;
                     //_\end_source
                     
                     //_\source ./warpv.tlv 1282   // Instantiated from warp-v_5-stage.tlv, 11 as: m4+riscv_csr(m4_echo(['m4_csr_']csr['_args']))
                        //--------------
                        // CSR TIME
                        //--------------
                        //_@0
                           assign FETCH_Instr_is_csr_time_a0 = FETCH_Instr_raw_a0[31:20] == 12'hC01;
                        //_@0
                           // CSR update. Counting on synthesis to optimize each bit, based on 32'b1.
                           
                           
                           // hw_wr_mask conditioned by hw_wr.
                           assign FETCH_Instr_csr_time_hw_wr_en_mask_a0[31:0] = {32{FETCH_Instr_csr_time_hw_wr_a0}} & FETCH_Instr_csr_time_hw_wr_mask_a0;
                           // The CSR value, updated by side-effect writes (if 1).
                           assign FETCH_Instr_upd_csr_time_a0[31:0] =
                                (FETCH_Instr_csr_time_hw_wr_en_mask_a0 & FETCH_Instr_csr_time_hw_wr_value_a0) | (! FETCH_Instr_csr_time_hw_wr_en_mask_a0 & FETCH_Instr_csr_time_a0);
                           // Next value of the CSR.
                           assign FETCH_Instr_csr_time_masked_wr_value_a0[31:0] =
                                FETCH_Instr_masked_csr_wr_value_a0[31:0] & 32'b1;
                           assign FETCH_Instr_csr_time_n1[31:0] =
                                FETCH_Instr_reset_a0 ? 32'b0 :
                                ((FETCH_Instr_is_csrrw_instr_a0 || FETCH_Instr_is_csrrwi_instr_a0) && FETCH_Instr_is_csr_time_a0)
                                       ? FETCH_Instr_csr_time_masked_wr_value_a0 | (FETCH_Instr_upd_csr_time_a0 & ! 32'b1) :
                                ((FETCH_Instr_is_csrrs_instr_a0 || FETCH_Instr_is_csrrsi_instr_a0) && FETCH_Instr_is_csr_time_a0)
                                       ? FETCH_Instr_upd_csr_time_a0 |   FETCH_Instr_csr_time_masked_wr_value_a0 :
                                ((FETCH_Instr_is_csrrc_instr_a0 || FETCH_Instr_is_csrrci_instr_a0) && FETCH_Instr_is_csr_time_a0)
                                       ? FETCH_Instr_upd_csr_time_a0 & ~ FETCH_Instr_csr_time_masked_wr_value_a0 :
                                // retain
                                         FETCH_Instr_upd_csr_time_a0;
                     //_\end_source
                     
                     //_\source ./warpv.tlv 1282   // Instantiated from warp-v_5-stage.tlv, 11 as: m4+riscv_csr(m4_echo(['m4_csr_']csr['_args']))
                        //--------------
                        // CSR TIMEH
                        //--------------
                        //_@0
                           assign FETCH_Instr_is_csr_timeh_a0 = FETCH_Instr_raw_a0[31:20] == 12'hC81;
                        //_@0
                           // CSR update. Counting on synthesis to optimize each bit, based on 32'b1.
                           
                           
                           // hw_wr_mask conditioned by hw_wr.
                           assign FETCH_Instr_csr_timeh_hw_wr_en_mask_a0[31:0] = {32{FETCH_Instr_csr_timeh_hw_wr_a0}} & FETCH_Instr_csr_timeh_hw_wr_mask_a0;
                           // The CSR value, updated by side-effect writes (if 1).
                           assign FETCH_Instr_upd_csr_timeh_a0[31:0] =
                                (FETCH_Instr_csr_timeh_hw_wr_en_mask_a0 & FETCH_Instr_csr_timeh_hw_wr_value_a0) | (! FETCH_Instr_csr_timeh_hw_wr_en_mask_a0 & FETCH_Instr_csr_timeh_a0);
                           // Next value of the CSR.
                           assign FETCH_Instr_csr_timeh_masked_wr_value_a0[31:0] =
                                FETCH_Instr_masked_csr_wr_value_a0[31:0] & 32'b1;
                           assign FETCH_Instr_csr_timeh_n1[31:0] =
                                FETCH_Instr_reset_a0 ? 32'b0 :
                                ((FETCH_Instr_is_csrrw_instr_a0 || FETCH_Instr_is_csrrwi_instr_a0) && FETCH_Instr_is_csr_timeh_a0)
                                       ? FETCH_Instr_csr_timeh_masked_wr_value_a0 | (FETCH_Instr_upd_csr_timeh_a0 & ! 32'b1) :
                                ((FETCH_Instr_is_csrrs_instr_a0 || FETCH_Instr_is_csrrsi_instr_a0) && FETCH_Instr_is_csr_timeh_a0)
                                       ? FETCH_Instr_upd_csr_timeh_a0 |   FETCH_Instr_csr_timeh_masked_wr_value_a0 :
                                ((FETCH_Instr_is_csrrc_instr_a0 || FETCH_Instr_is_csrrci_instr_a0) && FETCH_Instr_is_csr_timeh_a0)
                                       ? FETCH_Instr_upd_csr_timeh_a0 & ~ FETCH_Instr_csr_timeh_masked_wr_value_a0 :
                                // retain
                                         FETCH_Instr_upd_csr_timeh_a0;
                     //_\end_source
                     
                     //_\source ./warpv.tlv 1282   // Instantiated from warp-v_5-stage.tlv, 11 as: m4+riscv_csr(m4_echo(['m4_csr_']csr['_args']))
                        //--------------
                        // CSR INSTRET
                        //--------------
                        //_@0
                           assign FETCH_Instr_is_csr_instret_a0 = FETCH_Instr_raw_a0[31:20] == 12'hC02;
                        //_@0
                           // CSR update. Counting on synthesis to optimize each bit, based on 32'b1.
                           
                           
                           // hw_wr_mask conditioned by hw_wr.
                           assign FETCH_Instr_csr_instret_hw_wr_en_mask_a0[31:0] = {32{FETCH_Instr_csr_instret_hw_wr_a0}} & FETCH_Instr_csr_instret_hw_wr_mask_a0;
                           // The CSR value, updated by side-effect writes (if 1).
                           assign FETCH_Instr_upd_csr_instret_a0[31:0] =
                                (FETCH_Instr_csr_instret_hw_wr_en_mask_a0 & FETCH_Instr_csr_instret_hw_wr_value_a0) | (! FETCH_Instr_csr_instret_hw_wr_en_mask_a0 & FETCH_Instr_csr_instret_a0);
                           // Next value of the CSR.
                           assign FETCH_Instr_csr_instret_masked_wr_value_a0[31:0] =
                                FETCH_Instr_masked_csr_wr_value_a0[31:0] & 32'b1;
                           assign FETCH_Instr_csr_instret_n1[31:0] =
                                FETCH_Instr_reset_a0 ? 32'b0 :
                                ((FETCH_Instr_is_csrrw_instr_a0 || FETCH_Instr_is_csrrwi_instr_a0) && FETCH_Instr_is_csr_instret_a0)
                                       ? FETCH_Instr_csr_instret_masked_wr_value_a0 | (FETCH_Instr_upd_csr_instret_a0 & ! 32'b1) :
                                ((FETCH_Instr_is_csrrs_instr_a0 || FETCH_Instr_is_csrrsi_instr_a0) && FETCH_Instr_is_csr_instret_a0)
                                       ? FETCH_Instr_upd_csr_instret_a0 |   FETCH_Instr_csr_instret_masked_wr_value_a0 :
                                ((FETCH_Instr_is_csrrc_instr_a0 || FETCH_Instr_is_csrrci_instr_a0) && FETCH_Instr_is_csr_instret_a0)
                                       ? FETCH_Instr_upd_csr_instret_a0 & ~ FETCH_Instr_csr_instret_masked_wr_value_a0 :
                                // retain
                                         FETCH_Instr_upd_csr_instret_a0;
                     //_\end_source
                     
                     //_\source ./warpv.tlv 1282   // Instantiated from warp-v_5-stage.tlv, 11 as: m4+riscv_csr(m4_echo(['m4_csr_']csr['_args']))
                        //--------------
                        // CSR INSTRETH
                        //--------------
                        //_@0
                           assign FETCH_Instr_is_csr_instreth_a0 = FETCH_Instr_raw_a0[31:20] == 12'hC82;
                        //_@0
                           // CSR update. Counting on synthesis to optimize each bit, based on 32'b1.
                           
                           
                           // hw_wr_mask conditioned by hw_wr.
                           assign FETCH_Instr_csr_instreth_hw_wr_en_mask_a0[31:0] = {32{FETCH_Instr_csr_instreth_hw_wr_a0}} & FETCH_Instr_csr_instreth_hw_wr_mask_a0;
                           // The CSR value, updated by side-effect writes (if 1).
                           assign FETCH_Instr_upd_csr_instreth_a0[31:0] =
                                (FETCH_Instr_csr_instreth_hw_wr_en_mask_a0 & FETCH_Instr_csr_instreth_hw_wr_value_a0) | (! FETCH_Instr_csr_instreth_hw_wr_en_mask_a0 & FETCH_Instr_csr_instreth_a0);
                           // Next value of the CSR.
                           assign FETCH_Instr_csr_instreth_masked_wr_value_a0[31:0] =
                                FETCH_Instr_masked_csr_wr_value_a0[31:0] & 32'b1;
                           assign FETCH_Instr_csr_instreth_n1[31:0] =
                                FETCH_Instr_reset_a0 ? 32'b0 :
                                ((FETCH_Instr_is_csrrw_instr_a0 || FETCH_Instr_is_csrrwi_instr_a0) && FETCH_Instr_is_csr_instreth_a0)
                                       ? FETCH_Instr_csr_instreth_masked_wr_value_a0 | (FETCH_Instr_upd_csr_instreth_a0 & ! 32'b1) :
                                ((FETCH_Instr_is_csrrs_instr_a0 || FETCH_Instr_is_csrrsi_instr_a0) && FETCH_Instr_is_csr_instreth_a0)
                                       ? FETCH_Instr_upd_csr_instreth_a0 |   FETCH_Instr_csr_instreth_masked_wr_value_a0 :
                                ((FETCH_Instr_is_csrrc_instr_a0 || FETCH_Instr_is_csrrci_instr_a0) && FETCH_Instr_is_csr_instreth_a0)
                                       ? FETCH_Instr_upd_csr_instreth_a0 & ~ FETCH_Instr_csr_instreth_masked_wr_value_a0 :
                                // retain
                                         FETCH_Instr_upd_csr_instreth_a0;
                     //_\end_source
                     
                  //_\end_source
                  //_@0
                     //_\source ./warpv.tlv 1317   // Instantiated from warp-v_5-stage.tlv, 1529 as: m4+riscv_csr_logic()
                        
                        // CSR write value for CSR write instructions.
                        assign FETCH_Instr_masked_csr_wr_value_a0[31:0] = FETCH_Instr_raw_funct3_a0[2] ? {27'b0, FETCH_Instr_raw_rs1_a0} : L1b_FETCH_Instr_Src[1].L1_reg_value_a0;
                        
                     
                        // Counter CSR
                        //
                        
                        // Count within time unit. This is not reset on writes to time CSR, so time CSR is only accurate to time unit.
                        assign FETCH_Instr_RemainingCyclesWithinTimeUnit_n1[30-1:0] =
                             (FETCH_Instr_reset_a0 || FETCH_Instr_time_unit_expires_a0) ?
                                    30'd999999999 :
                                    FETCH_Instr_RemainingCyclesWithinTimeUnit_a0 - 30'b1;
                        assign FETCH_Instr_time_unit_expires_a0 = !( | FETCH_Instr_RemainingCyclesWithinTimeUnit_a0);  // reaches zero
                        
                        assign FETCH_Instr_full_csr_cycle_hw_wr_value_a0[63:0]   = {FETCH_Instr_csr_cycleh_a0,   FETCH_Instr_csr_cycle_a0  } + 64'b1;
                        assign FETCH_Instr_full_csr_time_hw_wr_value_a0[63:0]    = {FETCH_Instr_csr_timeh_a0,    FETCH_Instr_csr_time_a0   } + 64'b1;
                        assign FETCH_Instr_full_csr_instret_hw_wr_value_a0[63:0] = {FETCH_Instr_csr_instreth_a0, FETCH_Instr_csr_instret_a0} + 64'b1;
                     
                        // CSR write signals.
                        assign FETCH_Instr_csr_cycle_hw_wr_a0 = 1'b1;
                        assign FETCH_Instr_csr_cycle_hw_wr_mask_a0 = {32{1'b1}};
                        assign FETCH_Instr_csr_cycle_hw_wr_value_a0 = FETCH_Instr_full_csr_cycle_hw_wr_value_a0[31:0];
                        assign FETCH_Instr_csr_cycleh_hw_wr_a0 = 1'b1;
                        assign FETCH_Instr_csr_cycleh_hw_wr_mask_a0 = {32{1'b1}};
                        assign FETCH_Instr_csr_cycleh_hw_wr_value_a0 = FETCH_Instr_full_csr_cycle_hw_wr_value_a0[63:32];
                        assign FETCH_Instr_csr_time_hw_wr_a0 = FETCH_Instr_time_unit_expires_a0;
                        assign FETCH_Instr_csr_time_hw_wr_mask_a0 = {32{1'b1}};
                        assign FETCH_Instr_csr_time_hw_wr_value_a0 = FETCH_Instr_full_csr_time_hw_wr_value_a0[31:0];
                        assign FETCH_Instr_csr_timeh_hw_wr_a0 = FETCH_Instr_time_unit_expires_a0;
                        assign FETCH_Instr_csr_timeh_hw_wr_mask_a0 = {32{1'b1}};
                        assign FETCH_Instr_csr_timeh_hw_wr_value_a0 = FETCH_Instr_full_csr_time_hw_wr_value_a0[63:32];
                        assign FETCH_Instr_csr_instret_hw_wr_a0 = FETCH_Instr_commit_a0;
                        assign FETCH_Instr_csr_instret_hw_wr_mask_a0 = {32{1'b1}};
                        assign FETCH_Instr_csr_instret_hw_wr_value_a0 = FETCH_Instr_full_csr_instret_hw_wr_value_a0[31:0];
                        assign FETCH_Instr_csr_instreth_hw_wr_a0 = FETCH_Instr_commit_a0;
                        assign FETCH_Instr_csr_instreth_hw_wr_mask_a0 = {32{1'b1}};
                        assign FETCH_Instr_csr_instreth_hw_wr_value_a0 = FETCH_Instr_full_csr_instret_hw_wr_value_a0[63:32];
                        
                        
                        // For multicore CSRs:
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                        
                     //_\end_source
                     // CSR trap.
                     assign FETCH_Instr_is_csr_instr_a0 = FETCH_Instr_is_csrrw_instr_a0 ||
                                     FETCH_Instr_is_csrrs_instr_a0 ||
                                     FETCH_Instr_is_csrrc_instr_a0 ||
                                     FETCH_Instr_is_csrrwi_instr_a0 ||
                                     FETCH_Instr_is_csrrsi_instr_a0 ||
                                     FETCH_Instr_is_csrrci_instr_a0;
                     assign FETCH_Instr_valid_csr_a0 = FETCH_Instr_is_csr_instreth_a0 ? FETCH_Instr_csr_instreth_a0 : FETCH_Instr_is_csr_instret_a0 ? FETCH_Instr_csr_instret_a0 : FETCH_Instr_is_csr_timeh_a0 ? FETCH_Instr_csr_timeh_a0 : FETCH_Instr_is_csr_time_a0 ? FETCH_Instr_csr_time_a0 : FETCH_Instr_is_csr_cycleh_a0 ? FETCH_Instr_csr_cycleh_a0 : FETCH_Instr_is_csr_cycle_a0 ? FETCH_Instr_csr_cycle_a0 : 32'bx || FETCH_Instr_is_csr_instreth_a0;
                     assign FETCH_Instr_csr_trap_a0 = FETCH_Instr_is_csr_instr_a0 && FETCH_Instr_valid_csr_a0;
                     
                     // Memory inputs.
                     //_?$valid_exe
                        assign FETCH_Instr_unnatural_addr_trap_a0 = (FETCH_Instr_ld_st_word_a0 && (FETCH_Instr_addr_a0[1:0] != 2'b00)) || (FETCH_Instr_ld_st_half_a0 && FETCH_Instr_addr_a0[0]);
                     assign FETCH_Instr_ld_st_cond_a0 = FETCH_Instr_ld_st_a0 && FETCH_Instr_valid_exe_a0;
                     //_?$ld_st_cond
                        assign FETCH_Instr_addr_a0[31:0] = L1b_FETCH_Instr_Src[1].L1_reg_value_a0 + (FETCH_Instr_ld_a0 ? FETCH_Instr_raw_i_imm_a0 : FETCH_Instr_raw_s_imm_a0);
                        
                        // Hardware assumes natural alignment. Otherwise, trap, and handle in s/w (though no s/w provided).
                     assign FETCH_Instr_st_cond_a0 = FETCH_Instr_st_a0 && FETCH_Instr_valid_exe_a0;
                     //_?$st_cond
                        // Provide a value to store, naturally-aligned to memory, that will work regardless of the lower $addr bits.
                        assign FETCH_Instr_st_reg_value_a0[31:0] = L1b_FETCH_Instr_Src[2].L1_reg_value_a0;
                        assign FETCH_Instr_st_value_a0[31:0] =
                             FETCH_Instr_ld_st_word_a0 ? FETCH_Instr_st_reg_value_a0 :            // word
                             FETCH_Instr_ld_st_half_a0 ? {2{FETCH_Instr_st_reg_value_a0[15:0]}} : // half
                                           {4{FETCH_Instr_st_reg_value_a0[7:0]}};   // byte
                        assign FETCH_Instr_st_mask_a0[3:0] =
                             FETCH_Instr_ld_st_word_a0 ? 4'hf :                     // word
                             FETCH_Instr_ld_st_half_a0 ? (FETCH_Instr_addr_a0[1] ? 4'hc : 4'h3) : // half
                                           (4'h1 << FETCH_Instr_addr_a0[1:0]);      // byte
                     // Swizzle bytes for load result (assuming natural alignment).
                     //_?$returning_ld
                        //_/original_ld
                           // (Verilator didn't like indexing $ld_value by signal math, so we do these the long way.)
                           assign FETCH_Instr_OriginalLd_sign_bit_a0 =
                              ! FETCH_Instr_OriginalLd_raw_funct3_a0[2] && (  // Signed && ...
                                 FETCH_Instr_OriginalLd_ld_st_word_a0 ? FETCH_Instr_OriginalLd_ld_value_a0[31] :
                                 FETCH_Instr_OriginalLd_ld_st_half_a0 ? (FETCH_Instr_OriginalLd_addr_a0[1] ? FETCH_Instr_OriginalLd_ld_value_a0[31] : FETCH_Instr_OriginalLd_ld_value_a0[15]) :
                                               ((FETCH_Instr_OriginalLd_addr_a0[1:0] == 2'b00) ? FETCH_Instr_OriginalLd_ld_value_a0[7] :
                                                (FETCH_Instr_OriginalLd_addr_a0[1:0] == 2'b01) ? FETCH_Instr_OriginalLd_ld_value_a0[15] :
                                                (FETCH_Instr_OriginalLd_addr_a0[1:0] == 2'b10) ? FETCH_Instr_OriginalLd_ld_value_a0[23] :
                                                                        FETCH_Instr_OriginalLd_ld_value_a0[31]
                                               )
                              );
                           assign {FETCH_Instr_OriginalLd_ld_rslt_a0[31:0], FETCH_Instr_OriginalLd_ld_mask_a0[3:0]} =
                                FETCH_Instr_OriginalLd_ld_st_word_a0 ? {FETCH_Instr_OriginalLd_ld_value_a0, 4'b1111} :
                                FETCH_Instr_OriginalLd_ld_st_half_a0 ? {{16{FETCH_Instr_OriginalLd_sign_bit_a0}}, FETCH_Instr_OriginalLd_addr_a0[1] ? {FETCH_Instr_OriginalLd_ld_value_a0[31:16], 4'b1100} :
                                                                           {FETCH_Instr_OriginalLd_ld_value_a0[15:0] , 4'b0011}} :
                                              {{24{FETCH_Instr_OriginalLd_sign_bit_a0}}, (FETCH_Instr_OriginalLd_addr_a0[1:0] == 2'b00) ? {FETCH_Instr_OriginalLd_ld_value_a0[7:0]  , 4'b0001} :
                                                                (FETCH_Instr_OriginalLd_addr_a0[1:0] == 2'b01) ? {FETCH_Instr_OriginalLd_ld_value_a0[15:8] , 4'b0010} :
                                                                (FETCH_Instr_OriginalLd_addr_a0[1:0] == 2'b10) ? {FETCH_Instr_OriginalLd_ld_value_a0[23:16], 4'b0100} :
                                                                                        {FETCH_Instr_OriginalLd_ld_value_a0[31:24], 4'b1000}};
                           `BOGUS_USE(FETCH_Instr_OriginalLd_ld_mask_a0) // It's only for formal verification.
                     // ISA-specific trap conditions:
                     // I can't see in the spec which of these is to commit results. I've made choices that make riscv-formal happy.
                     assign FETCH_Instr_non_aborting_isa_trap_a0 = (FETCH_Instr_branch_a0 && FETCH_Instr_taken_a0 && FETCH_Instr_misaligned_pc_a0) ||
                                              (FETCH_Instr_jump_a0 && FETCH_Instr_misaligned_jump_target_a0) ||
                                              (FETCH_Instr_indirect_jump_a0 && FETCH_Instr_misaligned_indirect_jump_target_a0);
                     assign FETCH_Instr_aborting_isa_trap_a0 =     (FETCH_Instr_ld_st_a0 && FETCH_Instr_unnatural_addr_trap_a0) ||
                                              FETCH_Instr_csr_trap_a0;
                     
                  //_@0
                     // Mux the correct result.
                     //_\source ./warpv.tlv 1379   // Instantiated from warp-v_5-stage.tlv, 1593 as: m4+riscv_rslt_mux_expr()
                        assign FETCH_Instr_rslt_a0[31:0] =
                            FETCH_Instr_returning_ld_a0 ? FETCH_Instr_OriginalLd_ld_rslt_a0 :
                            32'b0 |
                            ({32{FETCH_Instr_is_lui_instr_a0}} & FETCH_Instr_lui_rslt_a0) |
                            ({32{FETCH_Instr_is_auipc_instr_a0}} & FETCH_Instr_auipc_rslt_a0) |
                            ({32{FETCH_Instr_is_jal_instr_a0}} & FETCH_Instr_jal_rslt_a0) |
                            ({32{FETCH_Instr_is_jalr_instr_a0}} & FETCH_Instr_jalr_rslt_a0) |
                            ({32{FETCH_Instr_is_lb_instr_a0}} & FETCH_Instr_lb_rslt_a0) |
                            ({32{FETCH_Instr_is_lh_instr_a0}} & FETCH_Instr_lh_rslt_a0) |
                            ({32{FETCH_Instr_is_lw_instr_a0}} & FETCH_Instr_lw_rslt_a0) |
                            ({32{FETCH_Instr_is_lbu_instr_a0}} & FETCH_Instr_lbu_rslt_a0) |
                            ({32{FETCH_Instr_is_lhu_instr_a0}} & FETCH_Instr_lhu_rslt_a0) |
                            ({32{FETCH_Instr_is_addi_instr_a0}} & FETCH_Instr_addi_rslt_a0) |
                            ({32{FETCH_Instr_is_slti_instr_a0}} & FETCH_Instr_slti_rslt_a0) |
                            ({32{FETCH_Instr_is_sltiu_instr_a0}} & FETCH_Instr_sltiu_rslt_a0) |
                            ({32{FETCH_Instr_is_xori_instr_a0}} & FETCH_Instr_xori_rslt_a0) |
                            ({32{FETCH_Instr_is_ori_instr_a0}} & FETCH_Instr_ori_rslt_a0) |
                            ({32{FETCH_Instr_is_andi_instr_a0}} & FETCH_Instr_andi_rslt_a0) |
                            ({32{FETCH_Instr_is_slli_instr_a0}} & FETCH_Instr_slli_rslt_a0) |
                            ({32{FETCH_Instr_is_srli_srai_instr_a0}} & FETCH_Instr_srli_srai_rslt_a0) |
                            ({32{FETCH_Instr_is_add_sub_instr_a0}} & FETCH_Instr_add_sub_rslt_a0) |
                            ({32{FETCH_Instr_is_sll_instr_a0}} & FETCH_Instr_sll_rslt_a0) |
                            ({32{FETCH_Instr_is_slt_instr_a0}} & FETCH_Instr_slt_rslt_a0) |
                            ({32{FETCH_Instr_is_sltu_instr_a0}} & FETCH_Instr_sltu_rslt_a0) |
                            ({32{FETCH_Instr_is_xor_instr_a0}} & FETCH_Instr_xor_rslt_a0) |
                            ({32{FETCH_Instr_is_srl_sra_instr_a0}} & FETCH_Instr_srl_sra_rslt_a0) |
                            ({32{FETCH_Instr_is_or_instr_a0}} & FETCH_Instr_or_rslt_a0) |
                            ({32{FETCH_Instr_is_and_instr_a0}} & FETCH_Instr_and_rslt_a0) |
                            ({32{FETCH_Instr_is_csrrw_instr_a0}} & FETCH_Instr_csrrw_rslt_a0) |
                            ({32{FETCH_Instr_is_csrrs_instr_a0}} & FETCH_Instr_csrrs_rslt_a0) |
                            ({32{FETCH_Instr_is_csrrc_instr_a0}} & FETCH_Instr_csrrc_rslt_a0) |
                            ({32{FETCH_Instr_is_csrrwi_instr_a0}} & FETCH_Instr_csrrwi_rslt_a0) |
                            ({32{FETCH_Instr_is_csrrsi_instr_a0}} & FETCH_Instr_csrrsi_rslt_a0) |
                            ({32{FETCH_Instr_is_csrrci_instr_a0}} & FETCH_Instr_csrrci_rslt_a0);
                     //_\end_source
                  
               //_\end_source
            
            //_@0
               
            //_@0
   
               // =======
               // Control
               // =======
   
               // Execute stage redirect conditions.
               assign FETCH_Instr_aborting_trap_a0 = FETCH_Instr_illegal_a0 || FETCH_Instr_aborting_isa_trap_a0;
               assign FETCH_Instr_non_aborting_trap_a0 = FETCH_Instr_non_aborting_isa_trap_a0;
               assign FETCH_Instr_mispred_branch_a0 = FETCH_Instr_branch_a0 && ! (FETCH_Instr_conditional_branch_a0 && (FETCH_Instr_taken_a0 == FETCH_Instr_pred_taken_a0));
               //_?$valid_decode_branch
                  assign FETCH_Instr_branch_redir_pc_a0[31:2] =
                     // If fallthrough predictor, branch mispred always redirects taken, otherwise PC+1 for not-taken.
                     
                     FETCH_Instr_branch_target_a0;
   
               assign FETCH_Instr_trap_target_a0[31:2] = 30'b0;  // TODO: What should this be?
               
               // Determine whether the instruction should commit it's result.
               //
               // Abort: Instruction triggers a condition causing a no-commit.
               // Commit: Ultimate decision to commit results of this instruction, considering aborts and
               //         prior-instruction redirects (good-path)
               //
               // Treatment of loads:
               //    Loads will commit. They write a garbage value and "pending" to the register file.
               //    Returning loads clobber an instruction. This instruction is $abort'ed (as is the
               //    returning load, since they are one in the same). Returning load must explicitly
               //    write results.
               //
               
               assign FETCH_Instr_abort_a0 = 1'b0 || FETCH_Instr_returning_ld_a0 || FETCH_Instr_replay_a0 || FETCH_Instr_aborting_trap_a0;  // Note that register bypass logic requires that abort conditions also redirect.
               // $commit = m4_valid_as_of(M4_NEXT_PC_STAGE + M4_MAX_REDIRECT_BUBBLES + 1), where +1 accounts for this
               // instruction's redirects. However, to meet timing, we consider this instruction separately, so,
               // commit if valid as of the latest redirect from prior instructions and not abort of this instruction.
               assign FETCH_Instr_commit_a0 = (! FETCH_Instr_reset_a0 && FETCH_Instr_next_good_path_mask_a0[(0 + 1) - 0]) && ! FETCH_Instr_abort_a0;
               
               // Conditions that commit results.
               assign FETCH_Instr_valid_dest_reg_valid_a0 = (FETCH_Instr_dest_reg_valid_a0 && FETCH_Instr_commit_a0) || FETCH_Instr_returning_ld_a0;
               assign FETCH_Instr_valid_ld_a0 = FETCH_Instr_ld_a0 && FETCH_Instr_commit_a0;
               assign FETCH_Instr_valid_st_a0 = FETCH_Instr_st_a0 && FETCH_Instr_commit_a0;
   
      //_\source ./warpv.tlv 1674   // Instantiated from warp-v_5-stage.tlv, 2059 as: m4+fixed_latency_fake_memory(/top, 0)
         // This macro assumes little-endian.
         
         //_|fetch
            //_/instr
               // ====
               // Load
               // ====
               //_@0
                  for (bank = 0; bank <= 4-1; bank++) begin : L1_FETCH_Instr_Bank //_/bank

                     // For $addr.
                     logic [31:0] L1_addr_a0;

                     // For $ld_value.
                     logic [(32 / 4) - 1 : 0] L1_ld_value_a0;

                     // For $spec_ld.
                     logic L1_spec_ld_a0;

                     // For $st_mask.
                     logic [3:0] L1_st_mask_a0;

                     // For $st_value.
                     logic [31:0] L1_st_value_a0;

                     // For $valid_st.
                     logic L1_valid_st_a0;

                     // For /mem$Value.
                     logic [(32 / 4) - 1 : 0] L1_Mem_Value_a0 [31:0];

                     assign {L1_addr_a0[31:0], L1_spec_ld_a0, L1_st_mask_a0[3:0], L1_st_value_a0[31:0], L1_valid_st_a0} = {FETCH_Instr_addr_a0, FETCH_Instr_spec_ld_a0, FETCH_Instr_st_mask_a0, FETCH_Instr_st_value_a0, FETCH_Instr_valid_st_a0}; // Find signal from outside of /bank.
                     //_/mem
                     //_?$spec_ld
                        assign L1_ld_value_a0[(32 / 4) - 1 : 0] = L1_Mem_Value_a0[L1_addr_a0[4 + 2 : 2]];
               
                     // Array writes are not currently permitted to use assignment
                     // syntax, so \always_comb is used, and this must be outside of
                     // when conditions, so we need to use if. <<1 because no <= support
                     // in this context. (This limitation will be lifted.)
      
                     // =====
                     // Store
                     // =====
      
                     /*SV_plus*/
                        always @ (posedge clk) begin
                           if (L1_valid_st_a0 && L1_st_mask_a0[bank])
                              L1_Mem_Value_a0[L1_addr_a0[4 + 2 : 2]][(32 / 4) - 1 : 0] <= L1_st_value_a0[(bank + 1) * (32 / 4) - 1: bank * (32 / 4)];
                        end
                  end
                  // Combine $ld_value per bank, assuming little-endian.
                  //$ld_value[M4_WORD_RANGE] = /bank[*]$ld_value;
                  // Unfortunately formal verification tools can't handle multiple packed dimensions produced by the expression above, so we
                  // build the concatination.
                  assign FETCH_Instr_ld_value_a0[31:0] = {L1_FETCH_Instr_Bank[3].L1_ld_value_a0, L1_FETCH_Instr_Bank[2].L1_ld_value_a0, L1_FETCH_Instr_Bank[1].L1_ld_value_a0, L1_FETCH_Instr_Bank[0].L1_ld_value_a0};
      
         // Return loads in |mem pipeline. We just hook up the |mem pipeline to the |fetch pipeline w/ the
         // right alignment.
         //_|mem
            //_/data
               //_@0
                  assign {MEM_Data_addr_a0[1:0], MEM_Data_dest_reg_a0[4:0], MEM_Data_ld_st_half_a0, MEM_Data_ld_st_word_a0, MEM_Data_ld_value_a0[31:0], MEM_Data_raw_funct3_a0[2], MEM_Data_valid_ld_a0} = {FETCH_Instr_addr_a0[1:0], FETCH_Instr_dest_reg_a0, FETCH_Instr_ld_st_half_a0, FETCH_Instr_ld_st_word_a0, FETCH_Instr_ld_value_a0, FETCH_Instr_raw_funct3_a0[2], FETCH_Instr_valid_ld_a0};
                  for (src = 1; src <= 2; src++) begin : L1_MEM_Data_Src //_/src

                     // For $dummy.
                     logic L1_dummy_a0,
                           L1_dummy_a1;

                     assign {L1_dummy_a0} = {L1b_FETCH_Instr_Src[src].L1_dummy_a0};
                  end
      //_\end_source
      //_|fetch
         //_/instr
            //_@0
               // =========
               // Reg Write
               // =========
   
               assign FETCH_Instr_reg_write_a0 = FETCH_Instr_reset_a0 ? 1'b0 : FETCH_Instr_valid_dest_reg_valid_a0;
               /*SV_plus*/
                  always @ (posedge clk) begin
                     if (FETCH_Instr_reg_write_a0)
                        FETCH_Instr_Regs_value_a0[FETCH_Instr_dest_reg_a0][31:0] <= FETCH_Instr_rslt_a0;
                  end
               
               // Write $pending along with $value, but coded differently because it must be reset.
               for (regs = 1; regs <= 31; regs++) begin : L1b_FETCH_Instr_Regs //_/regs
                  assign FETCH_Instr_Regs_pending_n1[regs] = ! FETCH_Instr_reset_a0 && (((regs == FETCH_Instr_dest_reg_a0) && FETCH_Instr_valid_dest_reg_valid_a0) ? FETCH_Instr_reg_wr_pending_a0 : FETCH_Instr_Regs_pending_a0[regs]);
               end
               
               
            //_@0
               `BOGUS_USE(L1_FETCH_Instr_OriginalLd_Src[2].L1_dummy_a0) // To pull $dummy through $ANY expressions, avoiding empty expressions.
   //_\end_source
   //_\source ./warpv.tlv 2082   // Instantiated from warp-v_5-stage.tlv, 12 as: m4+tb()
      //_|fetch
         //_/instr
            //_@0
               // Assert these to end simulation (before Makerchip cycle limit).
               assign FETCH_Instr_ReachedEnd_n1 = FETCH_Instr_reset_a0 ? 1'b0 : FETCH_Instr_ReachedEnd_a0 || FETCH_Instr_Pc_a0 == {30{1'b1}};
               assign FETCH_Instr_Reg4Became45_n1 = FETCH_Instr_reset_a0 ? 1'b0 : FETCH_Instr_Reg4Became45_a0 || (FETCH_Instr_ReachedEnd_a0 && FETCH_Instr_Regs_value_a0[4] == 32'd45);
               assign passed = ! reset && FETCH_Instr_ReachedEnd_a0 && FETCH_Instr_Reg4Became45_a0;
               assign failed = ! reset && (cyc_cnt > 200 || (! FETCH_Instr_reset_a3 && FETCH_Instr_commit_a6 && FETCH_Instr_illegal_a6));
   //_\end_source
endgenerate
//_\SV
   endmodule
